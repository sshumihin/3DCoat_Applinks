MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       sU�7x;�7x;�7x;ǩ���5x;�ƾ��x;�ƾ��wx;�ƾ���x;�7x:�mx;����2x;�����x;�����6x;�����6x;�Rich7x;�                PE  L ��OR        � !  �  `     ,4     �                         P         @                    � S   Lx <                            � <A  �� 8                           �Z @            � X                          .text   ��     �                   `.rdata  s�   �  �   �             @  @.data    F   �  &   j             @  �.reloc  rd   �  f   �             @  B                                                                                                                                                                                                                                                                                                                                                                                        V��舒 �N����*� �N$�2Z ��^���������������V��N$�����Z �N�W� ��^�o� ���������������j j j赲 �����U���   W���� ��u_��]�SVhx��M���Y �E�P�E�P�_$�} ��P�E�P�j^ ����P�/^ �M��wZ �M��oZ �M��gZ �G@    �x j S�E��Py �����Q  �E�P����Z P�M��Y �M�jj�E�Phtaoc�x ���M����Z ����MЋ@Q�@�Ѓ����M  ����M��@Q�@�С��j �@j��@�M�h��Q�С�����@�M��@8Q�wj���С���M��@Q�@�Ѓ��M��X �E�j	P��| ���M�P�*] �M��rY h���M��X h���M��X �E�P�E�P�E�P��p���P� ] ��P�E�P�] ����p����%Y �M��Y �M��Y �E�jP�
x ����t'�E�P�M��Y ���P�Qj�B8���ЍM��   ����M��@Q�@�С��j �@j��@�M�h��Q�ЍE�P�8 ����M��@Q�@�С���M��@Q�@�С��j �@j��@�M�h��Q�С����0�@�M��@8Qj���ЍM𡠴Q�@�@�С�����@j �@4j���С��j�@j�@0���С��j�@j�@0���С��j �@j�@0���С��j �@j�@0���С��j�@j�@0���С��j �@j
�@4���С��j�@j	�@0���С��j�@j�@0���С��j �@j�@0���С���M��@Q�@�С��j �@j��@�M�h��Q�С�����@�M��@8Qj���С���M��@Q�@�С�����@j �@0j���ЋM�V��o �M��u �M���V �M���V �_$�E�P���yW P�M��`V �M�jj�E�Phtaoc�ku ���M����V ����MЋ@Q�@�Ѓ���t3��  �M�j�wV��r �M��9u ����E�   �E�    �@�MЋ@Q�Ѓ��E�j j Pj�E�P���  P�E�P��膙 ����M��@Q�@�С���MЋ@Q�@�С���E�   �E�    �@�MЋ@Q�Ѓ��E�j j Pj�E�P���-  P�E�P���!� ����M��@Q�@�С���MЋ@Q�@�Ѓ��E�   �E�    h������h   ��@j ���   jh���h   �j j����P�E�P���4� ����E�   �E�    �@j ���   j j����P�E�P���ґ ����E�   �E�    �@j ���   j j����P�E�P��蠑 ����E�   �E�    �@j ���   j j����P�E�P���n� ����E�   �E�    �@j ���   j j����P�E�P���<� ����E�   �E�    j �@j ���   j����P�E�P���
� ���h���h   �j jh����E�
   �E�    �@h   ����   j j
����P�E�P���� ����E�	   �E�    �@j ���   j j	����P�E�P��萐 ����E�   �E�    �@j ���   j j����P�E�P���^� ����E�   �E�    �@j ���   j j����P�E�P���,� ����E�   �E�    �@�MЋ@Q�Ѓ��E�j j Pj�E�P���  P�E�P��虖 ����M��@Q�@�С���MЋ@Q�@�С�����E�   �E�    �@j ���   j j����P�E�P��蒏 h�  ���6� �   �E�P�Xq ����^[_��]�������������U����   SVW��3ۉ]��G@   �A  �E����   ����   H��  ����M��@Q�@�С��S�@j��@�M�h�Q�ЍE�P�� ����M��@Q�@���� h�h  h�   ���vN ��(��t��蘔  �ȍGPV�,�  _^�C[��]� �GP3�V��  _^�   [��]� �EP�E�P���E�   �]��m� 9]�  h�  ���� _^�   [��]� �� h�h�   j$����M ����t�@   ��X�X�X�X�3���WV���F  ����Mȋ@Q�@�С��j �@j��@�M�ht�Q�ЍE�P�� ����Mȋ@Q�@�С���M��@Q�@�С���� �@�M����   Qj�M�Q���Ћ�����I�E؋IP�ы���A�M؋@QV�С���M�@Q�@�С���M��@Q�@�С�����@j ���   j���Ѕ�tN����M��@Q�@�С��j �@j��@�M�h��Q�С�����@�M��@xQ�Mػ   �Ј]��u�E ��t����M��@Q�@�Ѓ��} �T  �Q  ������@��   �@dj�M��Ѝp�E�P�ƙRP�E���E��   �E�    ��  ������Qj�Rh��VW�M���j<��<���j P�G ����<���Pǅ<���<   ǅ@���    ǅD���    ǅH�������L���ǅT���    ǅX���   ǅ\���    �P���u4Ph����x����F  ��x���P�� �����x����@Q�@�Ѓ��EP�}�K ���@�@�M�Q�С��j �@j��@�M�h��Q�ЍE�P�v ����M��@Q�@�Ѓ�����M؋@Q�@�Ѓ�_^�   [��]� U���0W���@ t~V��l �E��E�P�O$�O P�M��N �M�jj�E�Phtaoc�m �MЋ��dN ����E�IP�I�у���^t����  �M��GP�g �M���l �E�P�l ��_��]���������������U���lW�E�P�E�P���E�   �E�    �|� �}� �\  V�M���L ����M܋@Q�@�С�����@�U܋��   Rj�U̍OR�Ћ�����I�E�IP�ы���A�M�@QV�С���M̋@Q�@�Ѓ��E�P�M���L �E�P�M��UP �M��MM ����M�@Q�@�С���M܋@Q�@�Ѓ��M�h���[L �E�P�M��/P �M��M �E�j P��k �����b  ����M�@S�@Q�С��j �@j��@�M�h��Q�ЍE�P�L ����M�@Q�@�Ѓ���j �߇ ����M�@Q�@�С��j �@j��@�M�h��Q�ЍE�jP�	 ������M�@Q�@���Ѓ� ��[��   ����M�@Q�@�С��j �@j��@�M�h�Q�ЍE�P� ����M�@Q�@���L� h�h�   h�   ���&H ��(��t	���H�  �3��OQV���؏  h�  ����� �M��K ^_��]� j j �E�P���E�   �E�    �� �M��K ^_��]� ���������������U���VW��j�wV�E�P�E�   �E�    艛 jV�E�P���E�   �E�    �m� jV�E�P���E�   �E�    聙 jV�E�P���E�   �E�    �� jV�E�P���E�   �E�    �� jV�E�P���E�   �E�    �͘ jV�E�P���E�   �E�    豘 jV�E�P���E�   �E�    蕘 j
V�E�P���E�
   �E�    �٘ j	V�E��E�	   �E�    P���]� jV�E�P���E�   �E�    �A� jV�E�P���E�   �E�    �%� jV�E�P���E�   �E�    �9� jV�E�P���E�   �E�    �� _^��]��������U���T  �H�3ŉE�Wj j�E ����u_�M�3���� ��]�V������PWǅ����(  �E ����   ������j�qE �����   ������QPǅ����$  �cE ��tt������P������h  P�� ������h  P�
� ���������P�@��u�+�/t��t������H��\uꍵ�����V�v� hp�V��� ����u.������PW��D ���F���W� �^3�_�M�3���� ��]ËM�^3͸   _��� ��]�������3���������������3������������������������������U��V��M�F   �F    � �9 u3�RQ���  ��^]� ��W�z�B��u�+�_RQ����  ��^]� ���������������U�졠�V�@��@V���u���j��@�u�@V�Ѓ���^]� ������������V��~r
�6��D ���F   �F    � ^�����������U��V��N$����|G �N��l ����~ �Et	V�D ����^]� �������U���EV�����t	V�hD ����^]� ��������������U��E�H�0����� Q�u�FC ��]��U��V�u�ƙ;�u 9Uu�E�H�0����� QV�C ��^]�3�^]��������������U�졠����@V���   W�u�U��uR�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]� �����������U��ESVW��������v���'�^������������;�v�����+��<;�v������G3ɉM��t���whjQQP�B �ȃ��E��tR�]��t�~r���ƅ�tSPQ�
� ���~r
�6��B ���E� ��~�^��r��_� ^[]� �<� ��U��E3Ʌ�t���wjQQP�B �ȃ���t��]� �� �U��S�]VW�{��M;���   +�9}B};�uG�9F��   �~�Fr�Qj ��� �  _��^[]� Q��j ��� �  _��^[]� �����   �F;�s$�v��W�����M��tj�{r��~r*��(��u�~��r�_�  ��^[]� _��^�  []� �օ�tW�PR��� ���~�~r��8 _��^[]� ���8 _��^[]� h���]� h���S� h���� ����������������U��S�]V���tW�N��r����;�rE��r���֋F�;�v1��r��u+�SV������^[]� �u��+�SV���q���^[]� W�}���w~�F;�s�v��W�`�����t_�~r*��(��u�~��r�_�  ��^[]� _��^�  []� �ƅ�tWSP�� ���~�~r��8 _��^[]� ���8 _��^[]� h���� ����������U��V�uV�Z� �����E�0t�@@�^]� �@H�^]� ���������������U��E�U��H]� ��������������U��E;Hu� ;Eu�]� 2�]� ��U�����U��uR�P�U�H;Ju� ;u���]� 2���]� �������������U��V��MW�~;�r~�U��+�;�w#�~�Nr�_� ��^]� ��_� ^]� ��tD�~r����+�S���+�tP�PS��� ���~�~[r��8 _��^]� ���8 _��^]� h����� �������U��V�u��� �u�������E��F   �F    � �: u3�QR���c�����^]� ��W�y��    �A��u�+�_QR���=�����^]� ������U��EV�u��u&j�F   �F    h4���� ������^]� PV�T�����^]� �������������U��V�u�e� �u�������E��F   �F    � �: u3�QR��������^]� ��W�y��    �A��u�+�_QR���}�����^]� �����̸������������̸(�����������̸h��������������������������������������������U��QV���F   �    �F    �F    �F    �F    �F(   �F    �F    �F,    �F$    �F     �F@   �F0    �F4    �FD    �F<    �F8    �FX   �FH    �FL    �F\    �FT    �FP    �Fp   �F`    �Fd    �Ft    �Fl    �Fh    ǆ�      �Fx    �F|    ǆ�       ǆ�       ǆ�       ǆ�      ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ǆ�      ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ���t�E��E�P�8; ���    �    �F    �F    �F    �F    �F��t�E��E�P��: ���F    �F    �F    �F,    �F$    �F     �F0��t�E��E�P�: ���F0    �F0    �F4    �FD    �F<    �F8    �FH��t�E��E�P�z: ���FH    �FH    �FL    �F\    �FT    �FP    �F`��t�E��E�P�:: ���F`    �F`    �Fd    �Ft    �Fl    �Fh    �Fx��t�E��E�P��9 ���Fx    �Fx    �F|    ǆ�       ǆ�       ǆ�       ���   ��t�E��E�P�9 ��ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ���   ��t�E��E�P�Y9 ��ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ��^��]����������U��QV���� ���   ��t�E��E�P��8 ��ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ���   ��t�E��E�P�8 ��ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       �Fx��t�E��E�P�78 ���Fx    �Fx    �F|    ǆ�       ǆ�       ǆ�       �F`��t�E��E�P��7 ���F`    �F`    �Fd    �Ft    �Fl    �Fh    �FH��t�E��E�P�7 ���FH    �FH    �FL    �F\    �FT    �FP    �F0��t�E��E�P�n7 ���F0    �F0    �F4    �FD    �F<    �F8    �F��t�E��E�P�.7 ���F    �F    �F    �F,    �F$    �F     ���t�E��E�P��6 ���    �    �F    �F    �F    �F    ^��]����������������U���  SVW��hG  �}��e# �O �����������u	_^[��]� �� �����8 ����M؋@Q�@�С���]�@�����   �M�Qj��p���Q���Ћ�����I�E��IP�ы���A�M��@QV�С����p����@Q�@�Ѓ��E�P�������8 �����P�� ����Z< ������O9 ����M��@Q�@�С���M؋@Q�@�ЋM�������P�{� P�� ����/< ������9 ����M��@Q�@�С���@�@j j��M�h��Q�Ѓ��E�P�� ����; ����M��@Q�@�Ѓ��������7 ����M؋@Q�@�С�����@�M؋��   Qj��p���Q���Ћ�����I�E��IP�ы���A�M��@QV�С����p����@Q�@�Ѓ��E�P������7 �����P�������; ������8 ����M��@Q�@�С���M؋@Q�@�Ѓ������h���7 �����P��������: ������7 ������6 ����M؋@Q�@�С�����@�M؋��   Qj��p���Q���Ћ�����I�E��IP�ы���A�M��@QV�С����p����@Q�@�Ѓ��E�P������6 �����P������: ������7 ����M��@Q�@�С���M؋@Q�@�Ѓ������h���6 �����P�������9 ������6 �E�P�� ����@7 P�:� ����M؋@Q�@�Ѓ��E�P�������7 P�� ����M؋@Q�@�Ѓ��E�P�������6 P��� ����M؋@Q�@������������PWɍ� ���P�E�P��(��������h���P������������� ����� ��������������E��M��M���h�����p�����x����i  ������   ���   �ЋMj P�E��u� ����M����   ���   �Ѕ��C  �RG ��h1D4ChCD4C�u��.� Pj j�����P���[: ����  ����M��@Q�@�С��j �@j��@�M�h��Q�Ѓ��E��u荍 �������P�E�P�5 PV�i  �����i  ����M؋@Q�@�С���M��@Q�@�С���M��@Q�@�С��j �@j��@�M�h��Q�Ѓ��E��u荍��������P�E�P�5 PV�i  ������  ����M؋@Q�@�С���@�M��@Q�С���M��@Q�@�С��j �@j��@�M�h��Q�С���u�@�����   j j����V����M�QP�E�P����b  PV�h  �����]  ����M؋@Q�@�С���M��@Q�@�С�����@j ���   j���Ѕ�t7�u衠����@��@V�С��j �@j��@h��V�Ѓ�����  ���j �@j���   ���Ѕ�t7�u衠����@��@V�С��j �@j��@h��V�Ѓ����  ���j �@j���   ����P�E�P����a  P�~� ����M؋@Q�@�ЋM���8 ����M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С��j �@j��@�M�h��Q�Ѓ�(�E�P��T���P�������2 P�E�P��p���P��f  ��P�E�P��f  P��� ����M؋@Q�@�С���@�@��p���Q�С����T����@Q�@�С���M��@Q�@�С���M��@Q�@�Ѓ�$�C ��h1D4ChCD4C�u��� Pj j�� ���P����6 ���V  ����M��@Q�@�С���M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�M�Q�С���M��@Q�@�С����$�@�u��@����V�С���M��@V�@Q�Ѓ����  ������d  �����P� ����M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С���@j �@j��M�h�Q�Ѓ�,�E�P�����P��T���h��P�z P�E�P��p���P�e  ��P�E�P�e  ����ЋA�M��@QR�С���M؋@Q�@�С����p����@Q�@�С����T����@Q�@�С���M��@Q�@�С���M��@Q�@�С����(�@�u��@����V�С��V�@�M��@Q�Ѓ����G  ����M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С��j �@j��@�M�h �Q�С����(�M�Q�0��T���P�l  P�E�P��p���P��c  ��P�E�P��c  ����ЋA�M��@QR�С���M؋@Q�@�С����p����@Q�@�С����T����@Q�@�С���@�@�M�Q�С���M��@Q�@�С����(�@�u��@����V�С���M��@V�@Q�Ћ������  �u����  ���j �@j���   �����F    �F    ���3����   �M����   ��H�����@����҅���  ��$    ��� ����M����   W���   �Ћ���؋��   �ˋR�]���=�  ��  ����������@Q�@�С��j �@j��@������h4�Q�С�������   �ˋ@x��P������P�����P�7b  P�q� ���������@Q�@�С���������@Q�@�Ѓ���<������������T����@Q�@�С��j �@j��@��T���hD�Q�С�������   �ˋ@x��P��T���P�� ���P�a  P�� ����� ����@Q�@�С���@�@��T���Q�Ѓ���H��� ��  ���h�  �@HS���   �Ѓ�������P�j  j�������j  ��������~
������3����E�    �O ���������}����
  �
��$    �I ������   �ϋ@��=�  ��  hF  h�  W����L  ����  j ���E�   �L �����$  h�  �u���p���P���M  �����p����@�@<�Ѕ��-  W�������i  �M�� �؉]���  �������������E����$    �d$ ������   �ˋ@��=)  ��   ����ˋ��   �@x�Ћ���ЋA��p����@xQ���Ѕ�ut���H ��d���Q��D���Qh���3�W�ȉE��B ��tI�]���I ��D���G;�d����M�I��@;�d���~�d���P��D���Ph���W���VB ��u]졠��ˋ��   �@(�Ћ؉E��� ����]�u���������������j �������8�`  �����p����@Q�@�Ћ}�������ϋ��   �@(�Ћ��E��������������? ��   ����M؋@Q�@�С��j �@j��@�M�hl�Q�С�������   �M؋@|Q�N �С���M؋@Q�@�С��j �@T�v �@�Ѓ����Z  �M�Q���u �������E��E��E��@�M��@HQh�  �M��ЋF �M����N �}� ��   ����   �������E�3�9~~T��    �F��������   �@x�Ћ�������   �E��Rx��ҋ���ЋAV�@x���Ћu���t8G;~|��}���E�F�E̅�x#jjjP����^  ��t�F�M̋U����}����}�K�c����]𡠴j �@Hh�  ��p  S�Ћ��j �IHh�  ��p  S�E��ы��h�  �IHS���   �E��ы��h�  �IHS���   �E��ы������؃�(�]�;�t(}+�QS�������f  �jj��+�PQ�������+^  3���~%�U���3�;B��������G�R���L��;�|ፅ<���P���RV  ��P����؋E쉝����;�t2}+�QP��<����h  ���P���jj+�PQ��<�����`  �����������0����@HQ�M��@8���������������������������������������������   ����h�����������Y��Y��Y��������Y��Y��Y���������8����������Y��Y��u��������Y��E��X��������X��������X��X��������������������X�8����E����������X��������������������������������Y��Y��Y��������Y��Y���0����������Y��������Y��Y�������������Y�������X��X��X��X��X�0�����8�����������X��}���8����������������������������������������������Y��������Y��Y��������Y��Y��Y���������L����������Y��Y��U�������������Y�������X��������X��������X��X���������������0����X�L�����������������X���������������������0�����x����Y��Y���L����������Y���p����Y��Y��Y���h����Y��������������Y��Y��������X��������X��������X��X��X��X��X�L����X��X������E���L�������������   �M̋�@����������}����
��$    �I �i��Q��f(��Y�����f(��Y�����Y�0����X��X�L���(��YE��X����������X�(��Y��X�(��Y�����Y�8���f�`��X�(��Y������Y��X��X��E��X�f�H�f�h�J�T���������;�t&��l���}+�PS�ia  �jj+�SP�
Y  �������u�3�3���~]�M�p������������<�u�A����D��A��D��A��D������A��D��A��D�������GT����;}�|��u�����M�@j ���   j�Ѕ���  ���j �@Hh'  �u����   �Ћ������q  ��h����E�;�t/��T���}+�PS�xb  �jj+�SP�i[  ��h����������E�������;�t)������}+�PS�O`  �jj+�SP��W  ��h����E���� ? W�3ɋ�3��U���0�����8�����@�����H�����P�����X�����`�����h�����p�����x����������������M����  ��X����I �����0����@DS�@,QR�ЋE􋍸������������<����   �~�x���f���~�����f�D��~�����f�D��~�`���f�D��~�h���f�D� �~�p���f�D�(�~�H����W�O�Rf���~�P���f�D��~�X���f�D��~�0����If���~�8���f�D��~�@���f�D��<��G�D����   �~�`���f���~�h���f�D��~�p���f�D��~�H���f�D��~�P���f�D� �~�X���f�D�(�~�0����O�If���~�8���f�D��~�@���f�D��G�<��D��������Ủ��M�A|���M�;M��\����]��u��u��u썅<���P�u����u��u��*  ��P���F����M�@j ���   j�Ѕ�t^��<����������@�������M����   G���   ��@�����;������]�M��a$ ��H��� t�~ ~S�u���79  ����M��@Q�@�ЍE�P��0 �E�P�E�    ��0 ����  ��h����!��������T����@Q�@�С��j �@j��@��T���hL�Q�С���M؋@Q�@�С��j �@j��@�M�hT�Q�С���M����   ��(�@x�Ѝ�T���QP�E�P�����P��R  ��P�� ���P��R  P��� ����� ����@Q�@�С��������@Q�@�С���M؋@Q�@�С����T����@Q�@�Ѓ� �o  �����p����@Q�@�С��j �@j��@��p���ht�Q�С���M؋@Q�@�С��j �@j��@�M�h��Q�С���M����   ��(�@x�Ћ�����I�E��IP�ы���A�M��@Q�M�Q�С�����@�M��@<�Ћ��j��Qj�VP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�Ѓ�����M��@�@<�Ћ��j��Qj���p���QP�BL�M��ЍE�P�P� ����M��@Q�@�С���M��@Q�@�С���M؋@Q�@�С����p����@Q�@�Ѓ���<������������M��@Q�@�Ѓ��E�P�>. ���E�    �E�P�+. ��3��[����M؋@Q�@�С��j �@j��@�M�h��Q�ЍE�P�� ����M؋@Q�@�Ѓ��������A ���   ������   �E����   P�у�������E�    � ������� �� ���� _��^[��]� ������������U�졠�S�@V�@dWj�M�ЍX�Ù�ȋ�;�u;�uh�h�  Q� �����3����j�@S�@hW�M��K3���~��7�MP��& F;�|�EP�}� ����M�@Q�@�Ѓ�_^[]� �������U�졠����@S�@V�M�WQ�С��j �@j��@�M�h��Q�С�����@j�@d�M��ЍX�Ù�ȋ�;�u;�uh�h�  Q� �����3����j�@S�@hW�M���K3���~�7�MP�& F;�|�EP�}� ����M��@Q�@�Ѓ�_^[��]� �����U���  ���S�@V�@W���M�Q�С��j �@j��@�M�ht�Q�С���M��@Q�@�С��j �@j��@�M�h��Q�ЋE��ء���ʋ@Q���   �M��M�SQ�]��Ћ�����I�E��IP�ы���A�M��@QV�С����@�@�M��@Q�С���MЋ@Q�@�С���MЋ@Q�M�Q�@�С�����@�MЋ@<�Ћ��j��Qj��M�QP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ��j��Qj��M�QP�BL�M��С���MЋ@Q�@�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�Ћ]������@S�@����V�С���M��@V�@Q�Ѓ��������u�E    �~ ��  �E    ������M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С��j �@j��@�M�h��Q�С����x����@Q�@�С��j �@j��@��x���h��Q�С����8����@Q�@�С����@�@j �@j���8���h��Q�ЋFE���������@���j0�@j ���   jj ���$Q�Ћ�����I������IP�ы���A������@QV�С���������@Q�@�ЋE��,�@Ej0j �@���j�@j ���   ���������$Q�Ћ�����I��(����IP�ы���A��(����@QV�С���������@Q�@�ЋE��,�@Ej0j � ���j�@j ���   ��������$Q�Ћ�����I��H����IP�ы���A��H���Q�@V�С��������@Q�@�С���M��@Q�@�С���M��@Q�@��8���Q�С����8�@�M��@<�Ћ��j��Qj���H���QP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ��j��Qj���x���QP�BL�M��С���M��@Q�@�С���M��@Q�M�Q�@�С�����@�M��@<�Ћ��j��Qj���(���QP�BL�M��С����h����@Q�@�С����h����@Q�@�M�Q�С�����@��h����@<�Ћ��j��Qj��M�QP�BL��h����С����X����@Q�@�С����X����@Q�@��h���Q�С�����@��X����@<�Ћ��j��Qj������QP�BL��X����С���MЋ@�@Q�С���MЋ@Q�@��X���Q�С�����@�MЋ@<�Ћ��j��Qj��M�QP�BL�M��С���M��@Q�@�M�Q�С���MЋ@Q�@�С����X����@Q�@�С����h����@Q�@�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С����H����@Q�@�С����(����@Q�@�С��������@Q�@�С����8����@Q�@�С����x����@Q�@�С���M��@Q�@�С���M��@Q�@�С����<�@S�@����V�С���M��@V�@Q�Ѓ��������E�u�E@�E;F�n��������x����@Q�@�С��j �@j��@��x���ht�Q�С���M��@Q�@�С��j �@j��@�M�h��Q�С���u��@�u����   �����Q�Ћ�����I�E��IP�ы���A�M��@QV�С����@�@������@Q�С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ���Qj�j��M�QP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ��j��Qj���x���QP�BL�M��С���M��@Q�@�M�Q�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С����x����@Q�@�С����S����@V�@�С���M��@V�@Q�Ѓ��������S����������M��@Q�@�Ѓ�_^[��]� ���������U���  ���S�@V�@�ٍM�WQ�]��С��j �@j��@�M�h��Q�С���M؋@Q�@�С��j �@j��@�M�h��Q�ЋE����@,�I�RP�E�P���   �Ћ�����I�EȋIP�ы���A�Mȋ@QV�С����@�@�M��@Q�С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ��j��Qj��M�QP�BL�M��С���M�@Q�@�С���M�@Q�@�M�Q�С�����@�M�@<�Ћ��j��Qj��M�QP�BL�M��С���M��@Q�@�С���Mȋ@Q�@�С���M؋@Q�@�С���M��@Q�@�С�����@�u�@����V�С���@�@�M�VQ�Ѓ���������u3�3��}�9]�a  �����(����@Q�@�С��j �@j��@��(���h��Q�С���������@Q�@�С��j �@j��@������h��Q�С���������@Q�@�С��j �@j��@������h��Q�С����h����@Q�@�С����@�@j �@j���h���h��Q�ЋF���<j0�D����j �@j���   j ���������$Q�Ћ�����I�������IP�ы���A�������@QV�С���������@Q�@�ЋE����@��,�\D����j0�@j ���   jj ���������$Q�Ћ�����I�������IP�ы���A�������@QV�С���������@Q�@�ЋE��,�@j0�����j �@j���   j ���������$Q�Ћ�����I��H����IP�ы���A��H���QV�@�С���������@Q�@�С����x����@Q�@�С����x����@Q�@��h���Q�С����8�@��x����@<�Ћ��j��Qj���H���QP�BL��x����С���������@Q�@�С���������@Q�@��x���Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������С���������@Q�@�С���������@Q�@������Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������С���������@Q�@�С���������@Q�@������Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������С���������@Q�@�С���������@Q�@������Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������С���M��@Q�@�С���M��@Q�@������Q�С�����@�M��@<�Ћ��j��Qj���(���QP�BL�M��С���M�@Q�@�M�Q�С���M��@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�С����x����@Q�@�С����H����@Q�@�С���������@Q�@�С���������@Q�@�С����h����@Q�@�С���������@Q�@�С���������@Q�@�С����(����@Q�@�С����<�@�u�@����V�С���M�@V�@Q�ЋM������������x����@Q�@�С��j �@j��@��x���h��Q�С���������@Q�@�С��j �@j��@������h��Q�С���@�������@Q�С��j �@j��@������h��Q�С��������@Q�@�С����@�@j �@j������h��Q�ЋE���@j0�D�(���j �@j���   j ����X����$Q�Ћ�����I�������IP�ы���A�������@QV�С����X����@Q�@�ЋE����@��,�\D� ���j0�@j jj ��������$Q���   �Ћ�����I��8����IP�ы���A��8����@QV�С��������@Q�@�ЋE��,�@j0�D����j �@j���   j ����8����$Q�Ћ�����I�������IP�ы���A�������@QV�С����8����@Q�@�С����h����@Q�@�С����h����@Q�@�����Q�С����8�@��h����@<�Ћ��j��Qj�������QP�BL��h����С����(����@Q�@�С����(����@Q�@��h���Q�С�����@��(����@<�Ћ��j��Qj�������QP�BL��(����С����H����@Q�@�С����H����@Q�@��(���Q�С�����@��H����@<�Ћ��j��Qj���8���QP�BL��H����С����H����@Q�@�С����H����@Q�@��H���Q�С�����@��H����@<�Ћ��j��Qj�������QP�BL��H����С����8����@Q�@�С����8����@Q�@��H���Q�С�����@��8����@<�Ћ��j��Qj�������QP�BL��8����С����X����@Q�@�С����X����@Q�@��8���Q�С�����@��X����@<�Ћ��j��Qj���x���QP�BL��X����С���M�@Q��X����@Q�С����X����@Q�@�С����8����@Q�@�С����H����@Q�@�С����H����@Q�@�С����(����@Q�@�С����h����@Q�@�С���������@Q�@�С����8����@Q�@�С���������@Q�@�С��������@Q�@�С���������@Q�@�С���������@Q�@�С����x����@Q�@�С����<�@�u�@����V�С���M�@V�@Q�ЋM����)������������@Q�@�С��j �@j��@�����h��Q�С���������@Q�@�С��j �@j��@������h��Q�С����(����@Q�@�С��j �@j��@��(���h��Q�С���������@Q�@�С����@�@j �@j�������h��Q�Ѓ��E�j0�<@�Ej �@j�D�@���j �@�����   ��x����$Q�Ћ�����I�������IP�ы���A�������@QV�С����x����@Q�@�ЋE����@��,�\D�8���j0�@j ���   jj ����h����$Q�Ћ�����I��X����IP�ы���A��X����@QV�С����h����@Q�@�ЋE��,�@j0�D�0����@���   j jj ����H����$Q�Ћ�����I�������IP�ы���A�������@QV�С����H����@Q�@�С����X����@Q�@�С����X����@Q�@������Q�С����8�@��X����@<�Ћ��j��Qj�������QP�BL��X����С���������@Q�@�С���������@Q�@��X���Q�С�����@�������@<�Ћ���Qj�j���(���QP�BL�������С���������@Q�@�С���������@Q�@������Q�С�����@�������@<�Ћ��j��Qj���X���QP�BL�������С���������@Q�@�С���������@Q�@������Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������С����h����@Q�@�С����h����@Q�@������Q�С�����@��h����@<�Ћ��j��Qj�������QP�BL��h����С��������@Q�@�С��������@Q�@��h���Q�С�����@������@<�Ћ��j��Qj������QP�BL������С���M�@Q�@�����Q�С��������@Q�@�С����h����@Q�@�С���������@Q�@�С���������@Q�@�С���@�@������Q�С����X����@Q�@�С���������@Q�@�С����X����@Q�@�С���������@Q�@�С���������@Q�@�С����(����@Q�@�С���������@Q�@�С��������@Q�@�С����<�@�u�@����V�С���M�@V�@Q�ЋM����?����u�F|�<���  ����M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С��j �@j��@�M�h��Q�С����x����@Q�@�С��j �@j��@��x���h��Q�С���������@Q�@�С����@�@j �@j�������h��Q�ЋE����<@�Fj0�D�X���j �@j���   j ����(����$Q�Ћ�����I�I������P�ы���A�������@QV�С����(����@Q�@�ЋE����@��,�\D�P���j0�@j ���   jj ��������$Q�Ћ�����I������IP�ы���A������@QV�С��������@Q�@�ЋE��,�@j0�D�H���j �@j���   j ���������$Q�Ћ�����I������IP�ы���A�����Q�@V�С���������@Q�@�С���Mȋ@Q�@�С���Mȋ@Q�@������Q�С����8�@�Mȋ@<�Ћ��j��Qj������QP�BL�M��С���M؋@Q�@�С���M؋@Q�@�M�Q�С�����@�M؋@<�Ћ��j��Qj���x���QP�BL�M��С���M��@Q�@�С���M��@Q�M�Q�@�С�����@�M��@<�Ћ��j��Qj������QP�BL�M��С���������@Q�@�С���������@Q�@�M�Q�С�����@�������@<�Ћ��j��Qj��M�QP�BL�������С��������@Q�@�С��������@Q�@������Q�С�����@������@<�Ћ��j��Qj�������QP�BL������С����8����@�@Q�С����8����@Q�@�����Q�С�����@��8����@<�Ћ��j��Qj��M�QP�BL��8����С���M�@Q�@��8���Q�С����8����@Q�@�С��������@Q�@�С���������@Q�@�С���M��@Q�@�С���M؋@Q�@�С���Mȋ@Q�@�С��������@Q�@�С��������@Q�@�С���������@Q�@�С���������@Q�@�С����x����@Q�@�С���M��@Q�@�С���M��@Q�@�С����<�@�u�@����V�С���M�@V�@Q�ЋM��������u�F|�}�<�C�}�;]����������x����@Q�@�С��j �@j��@��x���h��Q�С���M��@Q�@�С��j �@j��@�M�h��Q�ЋF,�����IRP������P���   �Ћ�����I�E��IP�ы���A�M��@QV�С����@�@�������@Q�С���M؋@Q�@�С���M؋@Q�@�M�Q�С�����@�M؋@<�Ћ��j��Qj��M�QP�BL�M��С���Mȋ@Q�@�С���Mȋ@Q�@�M�Q�С�����@�Mȋ@<�Ћ��j��Qj���x���QP�BL�M��С���M�@Q�@�M�Q�С���Mȋ@Q�@�С���M؋@Q�@�С���M��@Q�@�С���M��@Q�@�С����x����@Q�@�Ћ}��W������@��@V�С���M�@V�@Q�ЋM����x����M�W��������M�@Q�@�Ѓ�_^[��]� ��U���  ���S�@HV��p  Wj h�  �u���}��Ћ�����Q�M���   j j�E��ҋ���M�Rj ���   ��j��d����ҋ�����I�EЋIP��`����у�����  � ��  ��4����=�  ������P�q� ���z� P��4����.�  ��������  ����M��@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�P��4�����  ����M��@Q�@�С���M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С��j �@j��@�M�h��Q�Ѓ�,�E�P�E�P������P��4������  �����  P�E�P��x���P��'  ��P�E�P�'  ����ЋA�MЋ@QR�С���M��@Q�@�С����x����@Q�@�С���M��@Q�@�Ѓ� ���������  ����M��@Q�@�С���M��@Q�@�С�����@�u�@����V�С���MЋ@V�@Q�Ѓ���������u��������4����X�  ����M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С��j �@j��@�M�h��Q�С���M���   ��(�@x�Ћ�����I�E��IP�ы���A�M��@Q�M�Q�С�����@�M��@<�Ћ��j��Qj�VP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�Ѓ�����M��@�@<�Ћ��j��Qj��M�QP�BL�M��С���MЋ@Q�@�M�Q�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С�����@�u�@����V�С���MЋ@V�@Q�Ѓ����7����u��������u�uV�u�������ۋ]t�uȋ�SV�u�6��������h����@Q�@�С��j �@j��@��h���h��Q�С���M��@Q�@�С��j �@j��@�M�h��Q�Ћ���Ù�؋AR���   �M�SQ�]ȉU�Ћ�����I�E��IP�ы���A�M��@QW�С����@�@�M��@Q�С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�@<�M��Ћ��j��Qj��M�QP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ��j��Qj���h���QP�BL�M��С���MЋ@Q�@�M�Q�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С����h����@Q�@�С�����@�u�@����W�С���MЋ@W�@Q�Ћ}̃�������������$����@Q�@�E    �С��j �@j��@��$���h��Q�С����P����@Q�@�С��j �@j��@��P���h��Q��3ۃ�(�]9]��  ��I ��`��� �#  � �  ���   �����   ��������   �@x�Ћ���ЋA��P����@QR�С�����@��$����@xQ��P����Ѕ���  ����M��@Q�@�С��j �@j��@�M�h��Q�С����h����@Q�@�С��j �@j��@��h���h��Q�С���M��@Q�@�С���M��@Q�@��h���Q�С����4�@�M��@<�Ћ��j��Qj���P���QP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ���Qj�j��M�QP�BL�M��С���MЋ@Q�@�M�Q�С���M��@Q�@�С���M��@Q�@�С����h����@Q�@�С���M��@Q�@�С�����@�u�@����W�С���MЋ@W�@Q�Ћ}̃����n��������$����@Q�@��P���Q�Ѓ�����M��@Q�@�С��j �@j��@�M�h��Q�С���MЋ@Q�@�M�Q�С���M��@Q�@�ЋF|�� �<� �E    �|  �]�������������@Q�@�С��j �@j��@�����h��Q�С�����@�MЋ@<�Ћ��j��Qj������QP�BL�M��С��������@Q�@�ЋF4�O�A������IRP������P���   �Ћ�����I������IP�ы���A������@QW�С���������@Q�@�С���� �@�MЋ@<�Ћ��j��Qj������QP�BL�M��С��������@Q�@�Ѓ���d��� �%  �~\ �  ����M��@Q�@�С��j �@j��@�M�h��Q�С�����@�MЋ@<�Ћ��j��Qj��M�QP�BL�M��С���M��@Q�@�Ћ}̋FL�O�A������IRP��@���P���   �Ћ�����I��x����IP�ы���A��x����@QW�С����@����@Q�@�С���� �@�MЋ@<�Ћ��j��Qj���x���QP�BL�M��С����x����@Q�@�Ѓ��M�F|�U�}�A���M;�������ڡ���M��@Q�@�С��j �@j��@�M�h��Q�С�����@�MЋ@<�Ћ��j��Qj��M�QP�BL�M��С���M��@Q�@�С�����@�u�@����W�С���MЋ@W�@Q�Ћ}̃���������F|�M�C�M�];]�2�������M��@Q�@�С��j �@j��@�M�h��Q�С����x����@Q�@�С��j �@j��@��x���h��Q�С���u�@�uȋ��   ��@���Q�Ћ�����I�E��IP�ы���A�M��@QV�С����@�@��@����@Q�С���M��@Q�@�С���M��@Q�@��x���Q�С�����@�M��@<�Ћ���Qj�j��M�QP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ��j��Qj��M�QP�BL�M��С���MЋ@Q�@�M�Q�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С����x����@Q�@�С���M��@Q�@�Ћ]��S�������V�@�@�С���MЋ@V�@Q�Ѓ�������S���G��������P����@Q�@�С����$����@Q�@�С���MЋ@Q�@�Ѓ�_^[��]� ��U����   SV��W��8������  ����M̋@Q�@�С�����@�M̋��   Qj�M�Q�M�Ћ�����I�E�IP�ы���A�M�@QW�С���M��@Q�@�Ѓ��E�P��T������  ��T���P��8����:�  ��T����/�  ����M�@Q�@�С���M̋@Q�@�ЋM���E�P�^{ P��8�����  �M����  ����M�@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�P��8����m�  ����M�@Q�@�Ѓ��E�P��8�����  P�� ����M̋@Q�@�Ѓ��K�  ��h1D4ChCD4C�}��'� Pj j��8���P���T�  ��u3���  3ɉM9N��  �F������M܋@Q�@�С���M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С��j �@j��@�M�h��Q�С����,���   �ˋ@x�Ћ�����I�E�IP�ы���A�M�@Q�M�Q�С�����@�M�@<�Ћ��j��Qj�WP�BL�M��С���M��@Q�@�С���@�M��@Q�M�Q�С�����@�M��@<�Ћ��j��Qj��M�QP�BL�M��С���M܋@Q�@�M�Q�С���M��@Q�@�С���M�@Q�@�С���M��@Q�@�С���M��@Q�@�С�����@�u��@����W�С���M܋@W�@Q�Ѓ�������������p����@Q�@�С���@j �@j���p���h��Q�С���M܋@Q�@��p���Q�С����p����@Q�@�С���� �@�u��@����W�С���M܋@W�@Q�Ѓ����b���h�  S���u  ��tE������@���@W�С��j �@j��@h�W�Ѓ���h4  h@  S�u��u�,  h�  S���  ��tE������@���@W�С��j �@j��@h�W�Ѓ���h�	  hD  S�u��u��  �����`����@Q�@�С��j �@j��@��`���h�Q�С���M܋@Q�@��`���Q�С����`����@Q�@�С���� �@�u��@����W�С���M܋@W�@Q�Ѓ����$�������M��@Q�@�С��j �@j��@�M�h�Q�С���M܋@Q�@�M�Q�С���M��@Q�@�Ѓ� �u��������W�@�@�С���M܋@W�@Q�Ѓ�����������M̋@Q�@�С��j �@j��@�M�h,�Q�С���M܋@Q�@�M�Q�С���M̋@Q�@�С���� �@�u��@����W�С���M܋@W�@Q�Ѓ��������u�����������M܋@Q�@�ЋMA���M;N�?����M���  �   �E�P�D�  ����8����E�    �?�  _��^[��]� ����U���$�E�E�V�E�P�M��E�    �E�    �E�    �E�    �+ �Mj �E�P�E�P�	� �M���� ��tK����M܋��   Q�@X�Ћ�����t.����M���   �RT�ҋ���u�I|P�AV�Ѓ����3�����M܋��   Q� �Ѓ���^��]� ���������������U���$�E�E�V�E�P�M��E�    �E�    �E�    �E�    �[ �Mj �E�P�E�P�9� �M����� �����tU���   �M܋@HWQ�Ћ���}�IW�I���ы��W�IV�I�ы���E܋��   P�	�у���_^��]� �@�u�@V�С��j �Hj��Ih��V�ы���E܋��   P�	�у���^��]� ��������������U���$�E�E�V�E�P�M��E�    �E�    �E�    �E�    �[ �Mj �E�P�E�P�9� �M����� ��t����M܋��   Q�@8�Ѓ����3�����M܋��   Q� �Ѓ���^��]� ���������������U���$�E�E�    �E�S�E�P�M��E�    �E�    �E�    �E�    �  �Mj �E�P�E�P蒱 ��t����M܋��   Q�@�Ѓ���t��2ۍM�� ��[t����M܋��   Q�@<�Ѓ���E�E�E����]�M܋��   Q� ���E����]� ��������U���$�E�E�V�E�P�M��E�    �E�    �E�    �E�    ��� �Mj �E�P�E�P�ɰ �M����_ ��tS����M܋��   Q�@@���~ �u���f��~@���   f�F�~@�	�E�Pf�F�у���^��]� ����u���   W��	�E�P��F�F�у���^��]� ����U���$�E�E�V�E�P�M��E�    �E�    �E�    �E�    �� �Mj �E�P�E�P�� �M����  ��t"����M܋��   Q�@L�ЋM��P�[�  �
�Mj ���  ����E܋��   P�	�ыE��^��]� ��������������U���   ���S�@�ً@�M�VQ�С��j �@j��@�M�h��Q�С���MЋ@Q�@�С���MЋ@Q�@�MQ�С���� �@�MЋ@<�Ћ��j��Qj��M�QP�BL�M��С���M��@Q�@�Ѓ���\����u���uP��������M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С��j �@j��@�M�h��Q�С��������@Q�@�С��j �@j��@�����h��Q�С����l����@��<���   j0j jj ���������$Q�Ћ�����I��8����IP�ы���A��8����@QV�С���������@Q�@�С����d����@��,���   j0j jj ��������$Q�Ћ�����I��H����IP�ы���A��H����@QV�С��������@Q�@�С����\����@��,���   j0j jj ����d����$Q�Ћ�����I��(����IP�ы���A��(����@QV�С����d����@Q�@�С���M��@Q�@�С���M��@Q�@��(���Q�С����8�@�M��@<�Ћ��j��Qj������QP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ��j��Qj���H���QP�BL�M��С����t����@Q�@�С����t����@Q�@�M�Q�С�����@��t����@<�Ћ��j��Qj��M�QP�BL��t����С���M��@Q�@�С���M��@Q�@��t���Q�С�����@�M��@<�Ћ��j��Qj���8���QP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ��j��Qj��M�QP�BL�M��С���MЋ@�@<�Ћ��j��Qj��M�QP�BL�M��С���M��@Q�@�С���M��@Q�@�С����t����@Q�@�С���M��@Q�@�С���M��@Q�@�С���@�@��(���Q�С����H����@Q�@�С����8����@Q�@�С��������@Q�@�С���M��@Q�@�С���M��@Q�@�С����,�@�u�@����V�С���MЋ@V�@Q�Ѓ����j���h�  �u���u��������  h�  P������P���������������  j j ������P�M���  �MP������P��X���P�k P�� ����X����s�  �M��k�  ����M��@Q�@�С��j �@j��@�M�h��Q�С���M��@Q�@�С��j �@j��@�M�h8�Q�С���M��@Q�@�С���M��@Q�@�M�Q�С����4�@�M��@<�Ћ��j��Qj��MQP�BL�M��С���M��@Q�@�С���M��@Q�@�M�Q�С�����@�M��@<�Ћ��j��Qj��M�QP�BL�M��С���MЋ@Q�@�M�Q�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�С��j �@j�h���M��@Q�Ѓ�,��d���P�������f�  ������I�E��IP�ы���A�M��@QV�С�����@�M��@<�Ћ��j��Qj��M�QP�BL�M��С���MЋ@�@<�Ћ��j��Qj��M�QP�BL�M��С���M��@Q�@�С����d����@Q�@�С���M��@Q�@�С�����@�u�@����V�С���@�MЋ@VQ�Ѓ����m������������  ���������  ����MЋ@Q�@�С���M�@Q�@�Ѓ�^[��]�$ ����������U��S�]3ɋ��   3���~zV��rb�s|��WW�WɁ�  �yI���A��+����    �o���f���oD��f��;�|�f��fo�fs�_f��fo�fs�f��f~�;�}�s|�@;�|���^[]� ������������U�졠���   �@V�u�@V�С��j �@j��@h��V�ЋE����
��  �$��� �����`����@Q�@�С��j �@j��@��`���h��Q�Ѓ���`���P���v  ��`����  �����P����@Q�@�С��j �@j��@��P���h��Q�Ѓ���P���P���)  ��P����M  ����M��@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�P����  �M��  ����M��@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�P���  �M���  ����M��@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�P���c  �M��  ����M��@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�P���"  �M��I  ����MЋ@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�P����  �M��  ����M��@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�P���  �M���   ����M��@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�P���_  �M��   �����p����@Q�@�С��j �@j��@��p���h�Q�Ѓ���p���P���  ��p����<����M��@Q�@�С��j �@j��@�M�h�Q�Ѓ��E�P����  �M𡠴Q�@�@�Ѓ�����M��@Q�@�С��j �@j��@�M�h�Q�С�����@�΋@<�Ћȡ��j��Pj��RL�E�PQ���ҋ���E��IP�I�у���^��]� �I �� ՚ "� c� �� � &� g� �� � 3� ������������U��E�V��������|�����v3�^]ËE�0�H����� QV�u�4�  ��^]���������������U��EV�W���ϋ������������|�����v_3�^]ËE�0�H����� QW�u���  ��_^]����������������  �A   �A   �A    �A    �A    �������U��EW���A�A�A�A �A(�A0�A8�A@�AH�AP�AX�~ f��~@f�A�~@�Ef�A�~ f�A�~@f�A �~@�Ef�A(�~ f�A0�~@f�A8�~@�Ef�A@�~ f�AH�~@f�AP�~@f�AX��]� ����������U�졠�V�@�u�@V�С��V�@�u�@�С�����@�΋@<�Ћ��j��Qj��u�RLP���ҋ�^]������������U�졠�V�@��@<�Ћ��j��Rj��u��P�BL�Ћ�^]� ��������������U��V�u�ƙ;�u 9Uu�E�H�0����� QV��  ��^]�3�^]��������������U��Q3�9A~V�u�2@�R;A|�^]� ���������������U��QV����t�E��E�P��  ���    �    �F    �F    �F    �F    ^��]��������U���VW�}���y
_3�^��]� S�]���  �N;ϋ�O�Ӄ~ �U�u:h@�h'  hx�h  @�K� ���=�� t
�=�� t�[_3�^��]� ��;��]  )^�N�$  �A��~�   +��N����E�F�ʙEыʉE������U��E��U��U;�u�;M�u�;M�|�;U�r��Ù;�|�9Er��E�NFȋ�N�E�@��E�    ��u�E�P�������RP�E�>  ������U�RQP�E�@  �����ȃ���������F���F�N��~?+���P��+EÍ�P���P�Gh �N��    P��+E��PQ�-h ���I  ��P��+E��P���+  ��~��    P��v��P��g ���N����F�  �FH�~@�F��ȋF�U��E�E�M;���   	;M���   �����E����;��D����E�;��9���;E�0���	;M�%����Ù9U�����;�������E�@��E�    ��u�E�P�E�����RP�E�g  ������M�Q�u�E�i  P�M����ȃ����������F���F�E�F�F;�}�N+���P��P���P��f ���} t9�N;�}��+���P�Fj ��P�x ���N��    P��j Q�px ���M��N[_�   ^��]� ���������U���S�]W����y
_3�[��]� V�u����  �O;ˋ�O�փ �U�u:h@�h'  hx�h  @�� ���=�� t
�=�� t�^_3�[��]� ��;���  )w�O�a  �A���   +��O������G�ʙ�ыȉu����ɉE����������U�E����U�;�u�;�u�;M�|�;U�r��u�ƙ;��s���	9E��h����U�O�WʉO�E�@��E�    ��u/�E�P����ȋ����������RP�E�>  �����u��U�RQP�E�@  �����ȃ����������G�@���G�O��~J+Í@��P��+Eƍ@��P�3�@��P��d �O�[��P��+E�@��PQ�d ���  �@��P��+E�@��P�v�g  ��~�[��P��w�I��P�wd ���G�@��ȉG�A  �GH�@�G��ȋG�U���E�E��M�;���   	;M��   �E�ы��M����ЋE������E�U�M�;�������E;������;E������	;M�������ƙ9U�����;��������E�@��E�    ��u0�E�P�E���ȋ����������RP�E�g  �����u��M�Q�u��E�i  P������ȃ�����I����G�@���G�E��G�G;�}%�O+Í@��P�[��P�3�@��P�#c ���} tA�O;�}��+��I�@��P�Gj ��P��t ���v��P�G�[j ��P�t ���} t[�WW�;�}%�G�R�ȋ�+ʅ�t� �@�@��Iu�G�[�ȅ�~��$    ��t��A�A��Nu�M��O^_�   [��]� ����U�졠����H�EV�WRP�E�P���   �Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]��������������U��V��W�~��y_3�^]� jjjW������t�N�E��_�   ^]� ������U��Q�E;�u	�   ]� }+�RP�   ]� jj+�PR����]� ����������U��E��V����   ^��]� S�]W��xB�~;�};�> t6�N��u:h@�h�  hx�h  @��� ���=�� t
�=�� t�_[3�^��]� ��;�|�������_[�   ^��]� �;ǋ�LЋ�+����U;���   V��~�N��    PQ��P�` ���N��~���F;���   ������V�ǋ})F+ȉN�N+���QR��+�R�g` �E�P�v�E�@��6�E��  �E�    �t����ȃ�����,����F)~_���F[�   ^��]� �F+�HǙ��@���O��E;�}#�E�N+��+�����WP��P��_ �E��;F}?�M�QP�6�E�@��E��  �E�    ������ȃ����������F���F�E�F�})~_[�   ^��]� �������U��E��W�����   _��]� SV�u��xB�_;�};�? t6�O��u:h@�h�  hx�h  @�� ���=�� t
�=�� t�^[3�_��]� ��;�|�������^[�   _��]� �;Ë�LЋ�+����U;���   W��~�O�v��P�RQ��P�^ ���_��[�ȋO�G;��  �Ù���W����O)w+މ_�]+ˍI��P�vR��+�R�j^ �E�P�w�E�@��7�E��  �E�    ������ȃ���������G)_�@^���G[�   _��]� �G+�HÙ��@���K��E;�}-�U�O+�+ލ[��P�2�@��P�v��P��] �E��;G}B�M�QP�7�E�@��E��  �E�    �/����ȃ����������G�@���G�E�G�])_^[�   _��]� ������������������������������������������U������V�P��FP�B�Ѓ��N$�{�  �N@�s�  �N\�k�  �u�ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       ǆ�       �Fx    �F|    ǆ�       ǆ�   �������   ���   �E�P���   ���   �9^  ���   �����   ��^��]����U���V�����   �ܹ  ���   �ѹ  ���   ����t?�u��M�Q���   P��]  ���   覹  ��ǆ�       ǆ�       ǆ�       ���   ��t'P�u�  ��ǆ�       ǆ�       ǆ�       �N\��  �N@��  �N$��  ����H�FP�A�Ѓ�^��]����U���  �H�3ŉE��ES��V�C ���W�@�}���   j j	���Љ���j �@j���   ���ЉC���j �@j���   ���ЉC���j �@j
���   ���ЉC����������@Q�@�С�����@���������   Qj������Q���Ћ�����I�������IP�ы���A�������@QV�С���������@Q�@�С���H�CP������P�A�С���������@Q�@�С���������@Q�@�С���������@Q�@�С����$�@���������   Qj������Q���Ћ�����I�������IP�ы���A�������@QV�С���������@Q�@�Ѓ�������P������裹  ������P�K$��  �������	�  ����������@Q�@�С���������@Q�@�Ѓ�������h����  ������P�K$�߼  ������费  ����������@Q�@�С�����@���������   Qj������Q���Ћ�����I�������IP�ы���A�������@QV�С���������@Q�@�Ѓ�������P������襸  ������P�K@��  ��������  ����������@Q�@�С���������@Q�@�Ѓ�������h,���  ������P�K@��  ������趸  j�������9d  ������P�K$�*�  ����ЋAj �@hh�   ������Q���С���������@Q�@�Ѓ�������j@jP�������m�  ��H��� ����@�@��  ������Q�С��j �@j��@������h��Q�С���������@Q�@�С��j �@j��@������h��Q�Ѓ�(������P�K$�\�  ������I�������IP�ы���A�������@Q������Q�С�����@�������@<�Ћ��j��Qj�VP�BL�������С���������@Q�@�С���������@Q�@������Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������Ѝ�����P�l ����������@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�Ѓ�3��  ������Q�С��j �@j��@������hh�Q�С���������@Q�@�С��j �@j��@������hl�Q�Ѓ�(������P�K$豶  ������I�������IP�ы���A�������@Q������Q�С�����@�������@<�Ћ��j��Qj�VP�BL�������С���������@Q�@�С���������@Q�@������Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������Ѝ�����P��j ����������@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�Ѓ�������j h�   P�������m�  �������r�  ������P��o ������6  ����������@Q�@�С��j �@j��@������h<�Q�С���������@Q�@�С��j �@j��@������h��Q�С���������@Q�@�С��j �@j��@������Q������Q�Ѓ�<������P������P������P������P������P������P����P�ki ����������@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�Ѓ�$�l ������P���a3  ������P���  �{ t-���   +��   ���Q���������t����   ���  ���	>  �k j h  ��l ���   �������@Ǆ�������������H�A��������������ne  �������@Ǆ�������������X����QP�J艌����ǅX������N �M�����_^3�[�] ��]� ���������V���   ����  �   ^�����������U���d  �H�3ŉE�SVW��j��T����]  �G\�����Q�ȉ�����褲  ���j�@������@d�Ѝp�ƙ�ȋڙ;�u!;�uhP�h  Q��  ���؉�X����3ۉ�X������j�@V�@hS�������j@jS��T������  ������ ����@�@��  ��|���Q�С��j �@j��@��|���h��Q�С����l����@Q�@�С��j �@j��@��l���h��Q�Ћ�������(��4���P謱  ������I��\����IP�ы���A��\����@Q��l���Q�С�����@��\����@<�Ћ��j��Qj�VP�BL��\����С����H����@Q�@�С����H����@Q�@��\���Q�С�����@��H����@<�Ћ��j��Qj���|���QP�BL��H����Ѝ�H���P��e �����H����@Q�@�С����\����@Q�@�С����4����@Q�@�С����l����@Q�@�С����|����@Q�@�Ѓ�3��?  ��l���Q�С��j �@j��@��l���hh�Q�С����|����@Q�@�С��j �@j��@��|���h��Q�Ѓ�(��4���P�O\��  ������I��H����IP�ы���A��H����@Q��|���Q�С�����@��H����@<�Ћ��j��Qj�VP�BL��H����С����\����@Q�@�С����\����@Q�@��H���Q�С�����@��\����@<�Ћ��j��Qj���l���QP�BL��\����Ѝ�\���P�-d �����\����@Q�@�С����H����@Q�@�С����4����@Q�@�С����|����@Q�@�С����l����@Q�@�Ћ�T������@��`����T  �8���ǅ����    �������6�΋�������P������P�~X  ����Ή������R��t�j���������j
��@ �Ј�����������������j h�   P��T����  j������Ph����n ������   ������@P���   ���������   ��  ������P������h��P��i �����|����@Q�@�С��j �@j��@������Q��|���Q�С���H���   �P��|���P�A�С����|����@Q�@�Ћ��   ��,Ǆ�       ��  j������Ph���n ����u"���   ���P������h��P�i �  j������Ph����m ����u"���   ���P������h��P��h �i  j������Ph���m ����u"���   ���P������h��P�h �-  j������Ph���em ����u1���   �A0�P�A(�P�A �P������h��P�\h ����  j������Ph��m ����u1���   �AH�P�A@�P�A8�P������h�P�h ���  j������Ph���l ����u1���   �A`�P�AX�P�AP�P������h�P��g ���O  j������Ph,��l ����u1���   �Ax�P�Ap�P�Ah�P������h0�P�{g ���  j������Ph@��9l ����uW������P������hH�P�Ag ��������j P��4����b������H���   ���P��4���P�A�Ѝ�4����qj������PhT���k ����uy������P������h\�P��f ��������j P��l����2b������H���   �   �P��l���P�A�Ѝ�l������Q�@�@�Ћ��   Ǆ�      ����T����@��`����������X���������P�������9�  ����T����[u  j�������.U  �G@�����Q�ȉ�������  ���j�@������@d�Ѝp�ƙ�ȋڙ;�u!;�uhP�hd  Q菥  ���؉������3ۉ��������j�@V�@hS�������j@jS�������3  ������ �����l����@Q�@�  �С��j �@j��@��l���h��Q�С����|����@Q�@�С��j �@j��@��|���h��Q�Ћ�������(��l���P��H���P��  P��|���P��\���P������P��4���P����P��] �����4����@Q�@�С����\����@Q�@�С����H����@Q�@�С����|����@Q�@�С����l����@Q�@�Ѓ�$3���  �С��j �@j��@��l���hh�Q�С����|����@Q�@�С��j �@j��@��|���h��Q�Ѓ�(��l���P��H���P�O@��  P��|���P��\���P������P��4���P����P��\ �����4����@Q�@�С����\����@Q�@�С����H����@Q�@�С����|����@Q�@�С����l����@Q�@�Ћ�����3ɋ@��$��������������  ��$    �������6�΋�������P������P�>Q  ����΋��R��t�j����j
�@ ���Ј�,�����,���������j h�   P�������vx  ���   +��   ���Q��������3����   3���X������$    �����|����@Q�@�С��j �@j��@������Q��|���Q�С�����   �@���@x��|����R�Ћ���؋I��I��|���P�у�F�_  ���   +��   ��X������Q��������C���   �X���;��S���������j������Phh���f �����  ���   i��   �   �P������hx�P��a ���������@�������6�΋�������P������P�O  ����Ή������R��t�j���������j
��@ �Ј�0�����0���������j h�   P��������v  �����l����@Q�@�С��j �@j��@������Q��l���Q�С���H���   �   �P��l���P�A�Ѝ�l����  �����������j	������Ph���e ������   �������@�������6�΋�������P������P�N  ����΋��R��t�j����j
�@ ���Ј�D�����D���������j h�   P��������u  �����\����@Q�@�С��j �@j��@������Q��\���Q�Ћ��������i��   �P���   ���   �P��\���P�B�Ѝ�\������Q�@�@�Ѓ� �������@�������`�����������D���P��D���蘟  ���������n  S�E^ �������  �����4����@Q�@�С��j �@j��@��4���h<�Q�С����l����@Q�@�С��j �@j��@��l���h��Q�С����|����@Q�@�С��j �@j��@��|���SQ�С����H����@Q�@�С����@�@��H����@Q��l���Q�С�����@��H����@<�Ћ��j��Qj���|���QP�BL��H����С����\����@Q�@�С����\����@Q�@��H���Q�С�����@��\����@<�Ћ��j��Qj���4���QP�BL��\����Ѝ�\���P� W �����\����@Q�@�С����H����@Q�@�С����|����@Q�@�С����l����@Q�@�С����4����@Q�@�Ѓ��   ���������@Q�@�Ћ��������@Ǆ�������������H�A��������������{S  �������@Ǆ������������H�A艄���������Pǅ�������< �����������@Q�@�Ћ�T������@ǄT�������T����H�A���P��������� ǅd���\�t0��p���������9u ��������������������������+ɉ������ t��d����k  ������ǅd������t ���t��P��t�j���V��  ����T����@ǄT������T����������QP�J艌P���ǅ�������; �M�����_^3�[�J ��]����������������U������QSVW��3ۋ��   ���   +�����������.  3��u���O P�3 ����u@hG  �m� �𡠴������   ���   ���   E���P�B|�ЋO j j V�0 VS����   VS���  � V��Su��  ���  VS���  jj���K� ���j ���   j�@���Ћ��   +��   �u����Q��������C���   u�;�sW���   �#����@�M�@Q�С��j �@j��@�M�h��Q�ЍE�P�S ����M�@Q�@�Ѓ�3�_^[��]�_^�   [��]�����U�졠���0�@TS�@Wj �u���Ћ�����u_[��]� V�E�P���w� �u���i��   �P���   �� �P�BHh�  �M��Ћ��   �^���    tI����P���   P�B8h�  �M��ЍCP�M���  ����MЋ@Q�@<h�  �M��ЍM��B�  �E�P���� �M���  _�   [��]� ��U�졠���H�@S�@V�ٍM�WQ�С��j �@j��@�M�h��Q�ЋE���   i��   ȉE������@�U�@xR���   �Ћ���؋I��I�E�P�у�����  ����u�@Tj	�@V�Ћ�����u	_^[��]� j �E�Ph�  �M��E�    �E�    �� P���mq �M��� ����M苀�   Q�@8�Ѓ���uFP�E�Ph�  �M��E�   �E�   躿 P���Bq �M��� ����M؋��   Q� �Ѓ��E�P��艃 ����u�P���   ��P�P�BHh�  �M��С���E�   �E�   �@�M؋��   QhT  �M��С���M؋��   Q� �Ћ��   ����1�    tK����P���   �P�B8h�  �M��ЍCP�M�軚  ����M̋@Q�@<h�  �M��ЍM���  �E�P���� �M��g�  ����M苀�   Q� �Ѓ�_^�   [��]� ���U�졠���H�@S�@V�ٍM�WQ�С��j �@j��@�M�h��Q�ЋE���   i��   ȉE������@�U�@xR���   �Ћ���؋I��I�E�P�у����F  ����}�@Tj�@W�Ћ�����u	_^[��]� j �E�Ph�  �M��E�    �E�    �Ž P���-o �M��ſ ����M苀�   Q�@8�Ѓ���uFP�E�Ph�  �M��E�   �E�   �z� P���o �M��z� ����M؋��   Q� �Ѓ��E�P���I� �M��   ���    tI����P���   P�B8h�  �M��ЍCP�M��ߘ  ����M̋@Q�@<h�  �M��ЍM��>�  �E�P���� �M�苾  ����M苀�   Q� �Ѓ�_^�   [��]� �������U�졠���H�@S�@V�ٍM�WQ�С��j �@j��@�M�h��Q�ЋE���   i��   ȉE������@�U�@xR���   �Ћ���؋I��I�E�P�у�����  ����u�@Tj�@V�Ћ�����u	_^[��]� j �E�Ph�  �M��E�    �E�    �� P���Mm �M��� ����M苀�   Q�@8�Ѓ���uFP�E�Ph�  �M��E�   �E�   蚻 P���"m �M�蚽 ����M؋��   Q� �Ѓ�j �E�Ph�  �M��E�   �E�   �S� P����l �M��S� ����M؋��   Q� �Ѓ��E�P���" �M��   ���    tI����P���   P�B8h�  �M��ЍCP�M�踖  ����M̋@Q�@<h�  �M��ЍM���  �E�P����~ �M��d�  ����M苀�   Q� �Ѓ�_^�   [��]� U���L���S�@V�@��M�WQ�u��С��j �@j��@�M�h��Q�Ћ]���i��   ���   �@���@x���   �U�R��Ћ���؋I��I�E�P�у�����  ����u�@Tj�@V�Ћ�����u	_^[��]� j �E�Ph�  �M��E�    �E�    �Ź P���-k �M��Ż ����M䋀�   Q�@8�Ѓ���uFP�E�Ph�  �M��E�   �E�   �z� P���k �M��z� ����Mԋ��   Q� �Ѓ��E�P���I} �M�j ���   �M����   �^��E�Z�Ph  �E�   �E��� ��P�j �M��� ����Mԋ��   Q� �Ћu������   ���    tK����P���   �P�B8h�  �M��ЍFP�M��z�  ����Mȋ@Q�@<h�  �M��ЍM��ٔ  �E�P���| �M��&�  ����M䋀�   Q� �Ѓ�_^�   [��]� ��U���  �H�3ŉE�SV�uW��3�j��l�����������@���ǅ����    ǅ����    ǅ����    ��t�����������|�����?  j@jV��l����Jj  ����@�@9�������  ��p���Q�С��S�@j��@��p���h��Q�С���������@Q�@�С��S�@j��@������h��Q�С����`����@Q�@�С��S�@j��@��`���VQ�С���������@Q�@�С����@�@�������@Q������Q�С�����@�������@<�Ћ��j��Qj���`���QP�BL�������С����L����@Q�@�С���@�@��L���Q������Q�С�����@��L����@<�Ћ��j��Qj���p���QP�BL��L����Ѝ�L���P�IH �����L����@Q�@�С���������@Q�@�С����`����@Q�@�С���������@Q�@�С����p����@Q�@�Ѓ��������  ������Q�С��j �@j��@������hh�Q�С���������@Q�@�С��j �@j��@������hl�Q�С����`����@Q�@�С��j �@j��@��`���VQ�С���������@Q�@�С����@�@�������@Q������Q�С�����@�������@<�Ћ��j��Qj���`���QP�BL�������С����L����@Q�@�С���@�@��L���Q������Q�С�����@��L����@<�Ћ��j��Qj�������QP�BL��L����Ѝ�L���P�zF �����L����@Q�@�С���������@Q�@�С����`����@Q�@�С���������@Q�@�С���������@Q�@�С����\����@�������@���Q������ǅD���    ǅ\���    �С��ˋ@�������@��`���Q�С��j �@Shx���`���Q�@�Ѝ�`���P��H �����`����@Q�@�Ћ�l�����8�@��x�����
  �������6�΋�������P������P�K:  ����Ή������R��t�j���������j
��@ �Ј�<�����<���������j h�   P��l����{a  j������Ph���P �����   ������P������h��P�K ����������@����a�  ������P�O\�  ��������  �O\蟑  ������P�������-�  ������P�O\���  �������ӎ  ��	  j������Ph���P �����#  �����`����@Q�@�Ћ�������������������;�t7�I �~r�6裋  ���������F   �F    � ��;�uҋ����������� ������ǅ����   ǅ����    ƅ���� u3���������Q��I �A��u�+�Q������P��������I��jj������P��T����n:  ������r���������  ��������P���ă��     �@   �@    �@ ��T�����F�@   �@    �  ���tPQ��*  ����I�Dt�    ��8���P�5  ����������@�~r�6�����(����@Q�@�С��j �@j��@��(���VQ�С����`����@Q�@��(���Q�С����(����@Q�@�Ћ��   +��   ���   ���Q���������� ǅ����    �t\3��������ȡ����`����@R�@x�Ѕ���   �N+�������������   ���Q���������9�����������r��N+���Q��������B�P����i  ������   �p+��   ���Q�鋇�   �������i��   ��8����P��`���P�F�Ћ��   +��   ���Q��������H���������������>  ������Pǅ��������' �����`����@Q�@�Ѓ��  j������Ph����L ����u7C���������   ����+ˉ�������P������h��P��G ���@  j������Ph���L ����u;��D������   �v�ȍAP�APQ������h��P�}G ��F��D�����  j������Ph���4L ����ut��\������   �4@��΍APQ������h��P�*G ���   ΍AP�APQ������h��P�G ���   ����\D��$��\����D�]  j������Ph���K �����?  ���������������������t���   ����+ϋD�t��������������������������;�t8�d$ �{r�3��  ���������C   �C    � ��;�uҋ�����������P�������������DA��jj������P��T����6  ��������A��������P���ă��     �@   �@    �@ ��T�����P�7  ��$���P�r1  ��t�����������@;�t6��~r�6�P�  ���������F   �F    � ��;�uҋ�����������+������É�������x�������*��������H���������  ����  �pu  ��3�������������ǅ����    �������������������������������������"  �   ��    �������j/P��P���P���g#  P��t����K=  ��P�����;  ��t����r����P��G H��������������P�������d  ��h��W��'  ����t*�r�?W�G H��������������P��������c  �������������@���   ��D����D$�D��D$�ȋ��$�R��������������x����������������������������������������H����$R�P��H��� ��ǅ����    �x  ������+���������+ϋ��������������������������I ������ ���   �S�Lp���������D�v ���   �������S�Lp���������D9������� ���   �������S�Lp���������D9�v���   �������S�Lp��������������� ���   ��������Lp���������D9�v���   ��������Lp���������D9������ ���   ��������Lp���������D9�v���   ��������Lp���������D9������������������@�� ��������;�H���������������r  ����������t'P讂  ��ǅ����    ǅ����    ǅ����    ��������t'P�}�  ��ǅ����    ǅ����    ǅ����    �������������+8  ������Pǅ�������-! ����������l����@��x���������l����P  �����\����@Q�@ǅ����   �Ћ�t�������l����@Ǆl�������l����H�A���h��������� ǅ|���\�t0������������9u ��������������������������+ɉ������ t��|����5O  ������ǅ|������t ���t��P��t�j���V�4�  ����l����@Ǆl������l����H�A艄h���������Pǅ�������� ����t>��������;�t)��~r
�6�Ӏ  ���F   �F    � ��;�u�S貀  ����������tA������;�t.�~r
�6莀  ���F   �F    � ��;�u؋�����V�g�  ���M�������_^3�[�N. ��]� ǅ����   ���)  �   �������������j/P������P���  P��t�����7  ��������t>������������P�<  ��������  ��ǅ����    ǅ����    ǅ����    ��x�����+�t�������������*��������3�������C  ��	��$    ����������t���j��[j ��P������ǅ����   ǅ����    ƅ���� �<����uI���������   ������C�������+�����P�A ���������������ыL�pH�D���   ���   ������j ������C�����h��P�lN  ����u9���������tJ���������   ������C�������+�����P�7A ���������������ыL�pH�D�������������r�������Z~  ��C;����������������������@��������������;�����w�������������t�������������   �{r���Ӌ��������������   ��+���������R������������m@ �NpH�D9������+˸���*�����������vQ��h��S�>   ����t<�{r�������S���   ������@ �Np������H���������D��������������������������������U����  �H�3ŉE�SV�uW��j�������h+  j@jV��������U  ��@��� ����������@Q�@��  �С��j �@j��@������h��Q�С���������@Q�@�С��j �@j��@������h��Q�С���������@Q�@�С��j �@j��@������VQ�С���������@Q�@�С����@�@�������@Q������Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������С���������@Q�@�С���������@Q�@������Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������Ѝ�����P��3 ����������@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�С���������@Q�@�Ѓ�3���  �С��j �@j��@������h��Q�Ѝ�����P�6 ����������@Q�@�Ћ��������@�������7  ������6�΋�������P������P��'  ����΋��R��t�j����j
�@ ���Ј�����������������j jcP�������5O  j������Ph���r> ����u���   �G|����+ȋ��   �D�h�  j������Ph���9> ����u"���   ���   ����+ȋ��   �D�l�D  j������Ph����= ����uo���   ���   @P���   �-[  ���   ����+ȋ��   �D�d    ���   ����+ȋ��   �D�h    ���   ����+ȋ��   �D�l    �  j������Ph���t= ������  �Gxǅ����   ������������8�����u3���������Q�A��u�+�Q������P�������7��jj������P��8����9(  ������r��������x  ��������Pǅ����    ǅ����    ǅ����    ���ă��     �@   �@    �@ ��8�����F�@   �@    �  ���tPQ�  ����I�Dt�    ������P�1#  ������+���������*��������N��@����   t#��t~3���   ���   ����+ЍF�D�d����   ����+ȋ��   �D�d������� .  �������-  ������Pǅ������� ���������@�������������������E  �w|3ɋƻ   ����jj j ���Q�v  �Ѓ�����   �N�����   �BW�I�@��@�� �@y���   ����������@Q�@�С��j �@j��@������h8�Q�Ѝ�����P�E/ ����������@Q�@�Ћ���������t>������������P��2  �������v  ��ǅ����    ǅ����    ǅ����    �������[,  ������Pǅ�������] ��3��  3ҋ��   3ɉ��   ������jj j ���Q�u  ����t#�V���x�HW�J�A��A���Iy��3����   ����������@Q�@�С��j �@j��@������hP�Q�����   ������P����P������P������P����P�. ����������@Q�@�С���������@Q�@�С���������@Q�@�Ћ��   +��   ����������������8ǅ����    ���  3ۍS �s���   3ɋDd@����jj j ���Q�mt  ���   j�Dp���   3ɋDd@����j j ���Q�At  ���   �Dt����������@Q�@�С��j �@j��@������h\�Q�Ћ��   ����Dd�I�RP������P���   �Ћ�����I��@�I������P�ы���A�������@QV�С���������@Q�@�С���������@Q�@�С���������@Q�@������Q�С�����@�������@<�Ћ��j��Qj�������QP�BL�������Ѝ�����P�,, ����������@Q�@�С���������@Q�@�С���������@Q�@�Ћ��   +��   ��������������������Fº    ��������;��[x�r������   �������@Ǆ�������������H�A���������@��� ǅ����\�t0��������4���9u ��(�����,���������������+ɉ��<��� t�������@  ��$���ǅ�������t ���t��P��t�j���V�r  ���������@Ǆ�������������P����QP�J艌����ǅP������R �M�����_^3�[�E  ��]� ��U���$  �H�3ŉE�SV��W��l����=! �����`�����t���PWɍ�����P�����P���������������P������ǅx���    ��t�����|����������������������������$�����,������������������������������L����@Q�@�С��j �@j��@��L���h��Q�Ѝ�L���P��, �����L����@Q�@�Ћ��   3ɉ�h������   +θ�����������������  3���d������    ��{ �   �}��tz����������@Q�@�С��j �@j��@�M�Q������Q�Ћ�`�����������P�	 ��\�������������@Q�@�Ѓ���\��� t��\���P�gb ���u��u��p ������t�������  ������   �A�d����@��D���Q�С��j �@j��@��D���VQ�С�������   ��D����@|Q���С����D����@Q�@�С��������@Q�@�С��j �@j��@�����h��Q�С���H�E�RP��$���P���   �Ћ�����I��T����IP�ы���A��T����@QV�С����$����@Q�@�С��������@Q�@�С��������@Q�@�����Q�С����@�@������@<�Ћ��j��Qj���T���QP�BL������Ѝ����P�,' ���������@Q�@�С����T����@Q�@�С��������@Q�@�С���������@Q�@�С��j �@j��@������h��Q�С���H�E�RP������P���   �Ћ�����I�������IP�ы���A�������@QV�С���������@Q�@�С����@�@������@Q�С��������@Q�@������Q�С�����@������@<�Ћ��j��Qj�������QP�BL������Ѝ����P��% ���������@Q�@�С���������@Q�@�С���������@Q�@�С��j �@Hh�  ���   W�Ћ��j �IH�����   h�  W��|����у�(��p����E�    �M����   3������$    �E� �t�T�L�D�+�x���+�x���+�x���+�x����������E��������~�����f��� ���������~� ���f�C�M�@�E��[;�|���l�����t�����|���3�9U���   ��x����@����$    ���   ��������\������d�������Y��Y�������Y��X������Y��X�����B�X���$����Y��X����������X�������Y�f�v��X���,����Y��X�������Y�f�n��X���4����Y��X�f�N�;U��.����M�; ��  �}� ��  W�Q�������������������������������������������������������������������������O� ������p������A  �}� ǅ|���    �;  3҉U��I �M􋛌   �D
�<@�D
�4@�D
�@�E��D�   �@�~�fօ<����~D�fօD����~D�fօL����~�fօT����~D�fօ\����~D�fօd����~�fօl����~D�fօt����~D�fօ|����~�fօ�����~D�fօ�����~D�fօ������<���������󥋵p������� �����|����ЋAD�������@0QSR�ЋU�C�� ��;]艝|�����l����U��������t���j V����X ���j ���   j�@����j h�  ���?X ����   �����d����@Q�@�С��j �@j��@��d���h��Q�С�������   �ϋ@x�Ћ�����I��(����IP�ы���A��(����@Q��d���Q�С�����@��(����@<�Ћ��j��Qj�VP�BL��(����Ѝ�(���P�! �����(����@Q�@�С����d����@Q�@�Ѓ��{ ��  �����<����@Q�@�С��j �@j��@��<���h��Q�Ћ��   ���   +ȉ�|������Q�����������u>��<���P������@��@V�С��V�@��|����@�Ѓ���W�  �  �  ��<���P������@��@V�С��V�@��|����@�Ѓ���W�b  ���   +��   ���Q���������   �p���;���  �E��   h)  �!� ����|�������  ����������IP�I�ѡ��j �@j��@������h �Q�С���H�ǙRP��|���P���   �Ћ�����I��4����IP�ы���A��4����@QV�С����|����@Q�@�С����L����@Q�@�С����L����@Q�@������Q�С����<�@��L����@<�Ћ��j��Qj���4���QP�BL��L����С����<����@Q��L���Q�@�С����L����@Q�@�С����4����@Q�@�С���������@Q�@�С�������   ��<����@|Q��|����Ћ�|����z� �U�3���8�����~ �؋M�9<�uV���I �U�F;�|苝l�����t�����3��LT �Ѕ�t!��    ����򋁈   �ʋ@(�ЋЅ�u�V��|���V���T ���j ���   j�@���Ћ��   }���<���P������@��@V�С��V�@W�@�Ѓ�����t�����  ���   +��   ��p����E��   ���Q��������G�p���;��j�����t��������<����@Q�@�Ѓ���`���j j j W���t�  ���j ���   j�@���Ѝ�����Ph�   ǅ����    ǅ����    ǅ����    ǅ����    ǅ����    ��������������  ������������   ��x���E쉅x���� ���   ���   ��d�����h���+θ���������������x�d���9�h���������   _^[�M�3��� ��]á����<����@Q�@�Ѓ�3�_^[�M�3�� ��]��3 �M�_^3�3�[� ��]�U��M�%R ��t!V��������   �ȋR(�҅�u��^]� 3�]� ����������U���VW���Q� �N ���EP�c�  P���� �M���  ����M�@@Q�@$W�С�����@j�@4h�  �M��С��j�@h�  �@4�M��С���u�@h�  �@8�M��С��j�@h�  �@4�M��С��j�@@�M�@(QW�ЋM��3��0Q ��t%�
��$    �I ��������   �ȋB(�Ѕ�u�MVW�Q ���j ���   j�@���ЍM��_�  ����M�@Q�@�Ѓ�_^��]� ���U���P�H�3ŉE��E�MSVW�E��Ej3��E�W�E�3�3�P�M��]��u��]��4  �ȉM����u2�u��M��A  �E��M���M�_�H�M�^�H[�M�3�� ��]� �E�E�+�QW�u��M��E�   �E�    �E� �����E�;���   ;���   ��+˸���*���������;u�uj�M��+  �u��]���<Å���   �F   �F    � �s�G@tPWV� ���
���    �G�F�G�F�G   �G    � �p;u�uj�M��*  �u��]���tW�F   �F    � �}�s�E�@tP�E�PV� ����E��E�    �E�F�E��F�E�   �E�    �E� ���}��u�r�u��K`  ���}��M�jGW�E�P��2  �ȉE���������PW�u��M��E�   �E�    �E� �x���E�P�M��\?  �}�r�u���_  ���M��E���E��A�EĉA���M�_^3�[�� ��]� ��U��j�h�d�    P��`SVW�H�3�P�E�d�    �e�3��}��E� �]��uЋ�@�L8��t��Pj ���!  ����   ��p�t0�6�u����P�E�P�  ���E����R��t�j����E�x�xr� �  �E�    ��H�t �D$��|��t�E܃��s�E��������u��L8�mG  �ЉU܅�t�����   ���}��E������uЋ�@�D     �D$    �}� u����H˅��  �Aǃy8 u�����A�I#���   �E�   �E�D��E�P����   h���M��  h�n�E�P�E$ �ʋE�@�HH�a���Rj�M�*  �E�N�u���@�L8��F  �#����M��PыB���z8 u�����B�Bu��
��E������]�}�����j j ��# ��th���M��  h�n�E�P�# h���M���  h�n�E�P�# ��@�L08��t��R�ËM�d�    Y_^[��]�����������U��U�: u3����V�p�@��u�+�^�MPR�qj �R,  �����]�����������U��Q�E(V�u��u�uD���̃��A�j�j �E,�A   �A    P� �F���E���̃��A�j�j �E�A   �A    P� ���V�D   ��D�}$r�u�\  ���}@�E$   �E     �E r�u,�p\  ����^��]�������U��EV�u;E(t@��MD�EP�$<  �E��t'�MQP�s����ȃ���@�D�E�    E��E;E(u��}$�ED�r�u��[  ���}@�E$   �E     �E r�u,��[  ����^]����U��V�uW�};�tn�Ƥ   ����H�FP�A�С��V�@�@�С���H�F�P�A�С���H�F�P�A�С���H��\���P�A�Ё��   ����\���;�u�_^]����������������U���E�uP�� 3Ƀ������]����U��S�]W�};��G  V�u����    ���V�H�G�P�A�ЋG��F��F�G�F�~Gf�F �~Gf�F(�~Gf�F0�~G$f�F8�~G,f�F@�~G4f�FH�~G<f�FP�~GDf�FX�~GLf�F`�~GTf�Fh�~G\f�Fp�~Gdf�Fx����H���   P�GlP�A�С���H���   P�G|P�A�Ћ��   ���   ����H���   P���   P�A�С���H���   P���   P�A�Ћ��   ���   ���   �O��(���   ;��������^_[]ËE_[]����������������U��M�E+�V���4�    VQ�u� � ���^]� ������U��Q�u�E�j P�u�u�u�  ����]� ������������U��Q�u�E�j P�u�u�u�  ����]� ������������U��Q�u�E�j P�u�u�u�u  ����]� ������������U��j�h�d�    P��SVW�H�3�P�E�d�    �e��u�u��E�    �}��I ��t��t���  O�}���   �u���E������M�d�    Y_^[��]Ëu�};�t���  ���   ;�u�j j �a �����U��j�h0�d�    PQSVW�H�3�P�E�d�    �e��E�    �u�}�]��$    ��tS���(  O�}��x�]���E������M�d�    Y_^[��]�j j �� ������U��j�hP�d�    P��SVW�H�3�P�E�d�    �e��u�u��E�    �]�}��;�t ��tW��� 	  ���   �u���   �}���E������ƋM�d�    Y_^[��]Ëu�};�t��$    ����  ���   ;�u�j j �2 ������U��j�hp�d�    PQSVW�H�3�P�E�d�    �e��E�    �]�u�}��$    ;�tWS�M�  ��x�]��x�}���E������ËM�d�    Y_^[��]�j j � ����������������U��j�h��d�    P��SVW�H�3�P�E�d�    �e��u�u��E�    �]�}��;���   ����   �F    �F    �F   �F    �~r�����  �s�G@tPWV�� ���
���    �G�F�G�F�G   �G    �r��  ���u���}�l������  ���u���}�V����E������ƋM�d�    Y_^[��]Ëu�};�t�]V���  ��;�u�j j �r ������U��Q�u�j �u�u�u�Y�������]���U��Q�u�j �u�u�u���������]���U��W�}��tV�u�   �^_]� ����U��� �E(V�uD�uj��E�j �E,P�M��E�   �E�    �E� �;���E���̃��A�j�j �E��A   �A    P� ����}�r�u��T  ���Ej��E�j �EP�M��E�   �E�    �E� �����E���̃��A�j�j �E��A   �A    P� ����}�r�u��,T  ���E�P����� ��@�}$�ED�r�u�T  ���}@�E$   �E     �E r�u,��S  ����^��]������������U��V�u�~r
�6�S  ���F   �F    � ^]� ���U���SVWj �M��� �=x�����]���u/W�M���� 9=x�u���@����x��M��7� �=x��M�	;ys�A�4���ub�3��y t��� ;xs
�@�4���uD��t�M����� _��^[��]��u�E�P�  �����t*�u��5������RV�a� ���M��� _��^[��]�h���M��z h8o�E�P� ���������U���SVWj �M��� �=������]���u/W�M���� 9=��u���@�������M��7� �=���M�	;ys�A�4���ub�3��y t��� ;xs
�@�4���uD��t�M����� _��^[��]��u�E�P�&  �����t*�u��5������RV�a� ���M��� _��^[��]�h���M��z h8o�E�P� ���������U��Q�} VW���E�    t����Gp���j �@�w���V�H�A�D9���G    �G    �H��(  ��@�����H�A��D9����W  �F�F�F�F�F�F �\��FL �FE �F$�F,�N�N�F(�F0�    �F �     �F0�     �F�     �F�     �F,�     �FP    �|��FH��_�F@    ^��]� ��U��Q�} VW���E�    t�0��F`���S�@j ����~�HW�A�D1���F    �F    �H��'  ��]�@���$���H�A��D1����P   3����   D������u����t����[t���M�y�Qr�	PRQ���=  _��^��]� ���VWjj ��j j���O  ������tj�`� ����3��F�F�F�F�F�F �~4�F$�F,�N�N�F(�F0�    �F _�     �F0�     �F�     �F�     �F,�     ��^��U��V�uW���G   �G    � �~s�F@tPVW�� ���
���    �F�G�F�G�F   �F    ��_� ^]� �������������U��EV���F�@   �@    �  ���t#PQ���������I�D��t�    ^]� ��^]� �U�졠�S�@V�@��WS�С���}�@S�@W�ЋG�C�G�C�G�C�~G f�C �~G(f�C(�~G0f�C0�~G8f�C8�~G@f�C@�~GHf�CH�~GPf�CP�~GXf�CX�~G`f�C`�~Ghf�Ch�~Gpf�Cp�~Gxf�Cx������   �@V�@�С��V�H���   P�A�С�����   �@V�@�С��V�H���   P�A�Ћ��   ���   ������   �@V�@�С���H���   VP�A�С�����   �@V�@�С��V�H���   P�A�Ћ��   ��<���   _^��[]� �����̡��V�@��@V��W��F �F(�F0�F8�F@�FH�FP�FX�F`�Fh�Fp�Fx����H���   P�A�С���H���   P�A�С���H���   P�A�С���H���   P�A�Ѓ���^����������U���Vj ����� �F    �F 3��F    �F f�F�F    �Ff�F �F$�F(�F,�F0�E��tPV�� ����^��]� �EP�M��E<�� h�n�E�P�E�4��� ��������U��V�uWV���� ����F�G�F�G�����_^]� U��� �H�3ŉE��US�: V���E�   �E�    �E� u3���p�@��u�+�WPR�M���	���E�}��0�x�E�CE�E��E�P��� �}��{����s_r�u��	K  ���M�^�����3�[��� ��]� ������������U��V�u���� �4���^]� �����U��V�uWV���� ����F�G�F�G��_^]� ������V��~P �\�t�V�FD9u�F8�N<��F��F,+ɉ�~L t���&  ���v4��t ���t��P��t�j���V�,J  ��^��������VW���G��O��@�D8�$��G��P�B��D:��G�����  �w��G����t ���t��P��t�j���V��I  ���G��@�D8���G��H�A�D9�_^�������V����t'�vP�  �6�I  ���    �F    �F    ^��������������̡��V�P�񍆴   P�B�С���H���   P�A�С���H���   P�A�С���H���   P�A�С��V�@�@�Ѓ�^�����������V��V�� �F,����t	P� ���F,    �F$��t	P�| ���F$    �F��t	P�e ���F    �F��t	P�N ���F    �F��t	P�7 ���F    �F��t	P�  ���F    ��^�8� ��� ����������̋	��t��P��t�j������������U��VW�}��;�tQ���t'�vP�#  �6��G  ���    �F    �F    ���G�F�G�F�    �G    �G    _��^]� +I��A   +I���   +I��!  �U��V�������Et	V�G  ����^]� ���������������U��VW�y���wp�@�D0����F��H�A��D1��N������F�V�@�D0���F��H�A�D1������ ���Et	W�G  ����_^]� ��U��V��V������ ���Et	V��F  ����^]� �����U��V�q��V�@R�D���B�H�A�D������ ���Et	V�F  ����^]� �������U��VW�y��w`���N���V����Z� ���Et	W�SF  ����_^]� ��������U��V��W�~4����t ���t��P��t�j���W�F  ���Et	V� F  ��_��^]� �����U��V��W�����  �~4����t ���t��P��t�j���W�E  ���Et	V�E  ��_��^]� ����������U���EV���P�t	V�xE  ����^]� ��������������U��V��F�`���~
�v� �
y�v�9E  ���v�� ���E�P�t	V�E  ����^]� ���������������U��V���7
 �Et	V��D  ����^]� ���������������U��jj j �u�D  ��]������������D  ����������̡��j �@Hh�  ���   Q�Ѓ��+I��   +I���H�   +I���X�   ����������������������U��E�у�u�zr��E�M�]� �zr�P�EP�E�P�u� ��]� �������������̍A������    D���������������U��V�uW�};�t)��~r
�6��C  ���F   �F    � ��;�u�_^]� ��U��� �H�3ŉE�S�ك{@ �  �{E ��   �j��P���u2�[�M�3��]� ��]ù   �E� W�f�E�E��CE�V�M��E�   �@ W��}��K@�E��P�E�}�C}�u�Cu��PV�CHP�R �� tHt��tT2��R�CE �M��U�u����E�C�+�t�sP��V�E�C�jP�Z  ��;�uƀ{E t��u�Vj�M��  �v�����}�_^r�u��B  ����[�M�3��� ��]ËM�3Ͱ[�p� ��]����������������U���8SW�}3ۉ]���tb9u^VjSSj�A  ������t7�M�   �	��u����
�A��u�AP�M������F    ����3��7^��t�M������_�   [��]����������������U���HSW�}3ۉ]�����   9u}VjSSj�A  ������tV�M�   �	��u����
�A��u�AP�M��'����E�P�F    �`��p� �~ f�F�~@��f�F�3��7^��t�M��G���_�   [��]������������̋A�8 t�A,� ��3����������������U��V�q+1������������������"""+�;�s3�;uBu��^]� �;uBu��^]� ����̃��   ������U��}�AE ���AL�A�A�A�A�A�A �A$�A,�Q�Q�A(�A0�    �A �U�     �A0�     �A�     �A�     �A,�     ��t�B�A�A�B�Q�Q �A,�A0�QP�|��AH�A@    ]� ��̍A�A�A�A�A�A �A$�A,�Q�Q�A(�A0�    �A �     �A0�     �A�     �A�     �A,�     ���������U��ES�]V���F8    �F<����   ��<��   �����   Wjj j S��>  ������tqS�uW�]� ���F<��N8u�F�8�F�8�F,��F<�u7��F�׉8�F Eщ�F0��+�ˉ�F�8 u�F�8�F�     �F,�8�N<_^[]� �[� �V��Wj �F0    �F    �F    �F  �F   �F    �F     �F$    �F(    �F,    �/  jj j j��=  ������tj�)� ����~0_^�_�F0    ^��������������U��j�h��d�    P��HSVW�H�3�P�E�d�    �e����}��Hσy �  �I<��t�S  �} u��@�D8ts�t80�6�u����P�EP�8������؋���R��t�j����E�    ��@�L88�;&  �E���uj j��H���%  ��ȋC�HHu*�E�������Hσy ue��M�d�    Y_^[��]� ��@�L88�-&  렋M��PыB���z8 u�����B�Bu�O+��E������}��j j � �A���y8 u�����A�I#�u2��M�d�    Y_^[��]� �E�   �E�D��E�P��th���M��&���h�n�E�P� ��th���M�����h�n�E�P� h���M������h�n�E�P�y ������������̋AP��tP�%� Y��U��j�h��d�    PQSVW�H�3�P�E�d�    �e����E�    ��@�|0 u%�D0t�L08��P4���uj j��H��M$  �E������M�d�    Y_^[��]ø�,��������������̋A �8 t�A0� ��3����������������U��j�h��d�    P��SVW�H�3�P�E�d�    �e���3��u�]��t*�����?wjVV��    P�:  �����u��u�� �E�    V�w�7���y����E�������G+����E��t	Q�;  �����G�E���G�7�M�d�    Y_^[��]� �u���:  ��j j ��  ���������������U��j�h�d�    P��SVW�H�3�P�E�d�    �e���3��}�u��t+���GwjWW��i��   P��9  �����}��u��� �E�    W�s�3��������E������K+���Q��������E���t�u�EP�sQ�B����3�:  ���E�i��   ��si��   ǉC�;�M�d�    Y_^[��]� �u���9  ��j j ��� �����U��j�h0�d�    P��SVW�H�3�P�E�d�    �e���3��u�}��t-��"""w jVV����+���P��8  �����u��u��� �E�    V�s�3��������E������K+��������������ʉM���tP�9  ���M����+ǍƉC����+��ƉC�3�M�d�    Y_^[��]� �u���8  ��j j ��� ��������������U��j�hP�d�    P��SVW�H�3�P�E�d�    �e���3��u�]��t)�����
wjVV�[��P��7  �����u��u��� �E�    V�w�7���*����E������O+����*��������ʉM���t�wP���9����7�8  ���M�[�ƉG�I�ƉG�7�M�d�    Y_^[��]� �u���7  ��j j ��� ����������������U��QV�q��+�W�}��;�sI+1S����?����+�;�r<+�������+�;�[s3�;�_B�^�U]������;�_B�^�U]����_^]� h����� ��������������U��S�YV�q��+ָ��Q��������W�}�;�sh+1���Q����������G+�;�rQ+���Q���������������G+�;�s3�;�_B�^[�E]�����;�_B�^[�E]�����_^[]� h���J� ���������������U��SVW��������_�w+���֋u�������;�s3+��������������ʸ"""+�;�r�1P���;���P���s���_^[]� h����� ��U��S�YV�q��+ָ���*��������W�}�;�sh+1����*��������򸪪�
+�;�rQ+����*�������������꿪��
+�;�s3�;�_B�^[�E]������;�_B�^[�E]�����_^[]� h���*� ���������������V�q�AD9u�A8�Q<��A��A,+҉^����������������V��W�z�rD�;�t�J�B8�B,� �B<�7�B�ʉ0�B,+΃�E_�^�����������V���F<t�F�0��4  ���F�     �F�     �F,�     �F�     �F �     �F0�     �f<��F8    ^��������U���V����t.�u��M�Q�vP�����6�z4  ���    �F    �F    ^��]���������������V����tP�A4  ���    �F    �F    ^��������̋AP��tP�T� Y��U��S�]V�����N+�;�v|��tpW�<���wy�F;�s3QW���]�����tR�u��S�v�{����~�~r5��8 _��^[]� ��u։~��r�_�  ��^[]� _��^�  []� ���8 _��^[]� h���� h���� ����������U��E���A�I��#�t!�E��E�   �E�D�P��u���M�u#�9��]� h���M�����h�n�E�P�� h���n���h�n�E�P��� h���V���h�n�E�P��� ��������U��E���A�I��#�t'�} u'�E��E�   �E�D�P��u���M�u,�B��]� j j �� h���M������h�n�E�P�u� h�������h�n�E�P�]� h������h�n�E�P�E� ���������V��W�~P u3�� �}����vP3Ʉ���D��*� 3Ƀ���E��F�F�F�F�F�F �FL �FE �F$�F,�N�N�F(�F0�    �F �     �F0�     �N���    �N_�    �N,�    �FP    �|��NH�F@    ^��������U���V��N�?�����uE��H�D1΃��y8 u�����A�I#�t!�E��E�   �E�D�P��u���M�u"�8^��]�h���M�����h�n�E�P�� h���l���h�n�E�P��� h���T���h�n�E�P��� ������U��A�U;�rLV�u+�;�B��yWr�	�}��;�B�P�u�P�8   ����u;�s	_���^]� 3�;���_^]� h���F� �������������U��M��u3�]ËUV�u��r��    �;u������s���t5�:u'���t*�B:Fu���t�B:Fu���t�B:Ft���^]�3�^]�U��E��tjxj P�<� ��]� ����̰�������������̸   �����������U��M�E��M �E��   ]� ����U��E+E9EBE]� ������������U��E]� ������U��U�M+�QR�u�[� �E��]� �U��AP�EP�� ��]� ��������U��V�uW�};�tS�Y�SP�~� �F��;�u�[_��^]� U��AP�EP�W� ��]� ��������U��V�uW�};�tS�Y�SP�+� �F��;�u�[_��^]� U��M�E�3�]� ���������������U��E]� ������U��U�M+�QR�u�k� �E��]� �U��Q�E�UVW���;�u-�w;�u&�u�E�PVQ�W�����M���G�E_�^��]� ;�t5�uP�wR������u���E�P�wV�����E�M�� �w_�^��]� �M_���^��]� �������U����U�EV�1�M�;�u;Au�E�q�^��]� ;�t2�qS��;�t$��W��I ������x�   ��x�;�u�U�M�_�Y[�E^���]� ����U��Q�US�]�M���u;Qw	��[��]� V�qW;�sj+�;�wd�   +���yr�	���tL�EV� PS��� ������t5�u�uW��������t
+�K�_�ȋE��xr� +���_^[��]� _^���[��]� �U���V���@�L08����   ��P��@�|0 u�L0<��t�������H�|1 ����tS�L18��P4���uE��H�D1΃��y8 u�����A�I#�t!�E��E�   �E�D�P��u3���M�uF�\�� ��u��������@�L08��t��P��^��]�h���M��N���h�n�E�P��� h���6���h�n�E�P��� h������h�n�E�P�� ����������������U��QSVW����@�t80�6�΋�u��P�E�P���������΋��R��t�j����j
�@ ���ЈE��u����u�u�u�   _^[��]� �������U��j�hp�d�    P��XSVW�H�3�P�E�d�    �e���u�3��}�~�~�u؋�@�L08��t��Pj���w�������   9}|�]��tv�E�E�E�    ��@�L08�%  �ȉM���u���A;Mu�F�V ��@�L08��  �'����]�E����E����   |����   ���}��E������E�  �FFu����H΅���   �Aǃy8 u�����A�I#���   �E�   �E�D��E�P����   h���M��D���h�n�E�P��� �F�V �E�@�E��@�L08�  �����M��PыB���z8 u�����B�Bu��>��E������u�}��+���j j �i� ��th���M�����h�n�E�P�I� h���M�����h�n�E�P�.� �M؋�@�L8��t��P�ƋM�d�    Y_^[��]� �������U��VW�u���A���������ϋR�҄�t_�F@    ^]� �Ή~@����_^]� ��� �������������U���SVW�������E�w0�G8�G<    �6�΋�u�P�EP���������΋��R��t�j����j �@ ���Ѓ8 �G@u4�G�O�����G#�t!�E��E�   �E�D�P��u"���M�u5�K�} t	W�� ��_^[��]� h���M��V���h�n�E�P��� h���>���h�n�E�P��� h���&���h�n�E�P�� ��������U��W���P uz�u�u�u�� ����teSVjP��������w4�6�΋�u�P�EP�����؃���ˋR�҄�t	�G@    �
�ω_@�6�������P^[��t�j�����_]� 3�_]� ���U��E����V�u��P�u�N�R�������HuG�D1΃��y8 u�����A�I#�tq��us�E����E�   �E�D�P�M���   �   3�9D18�   D��D1�L1#�t,��u/�E����E�   �E�D�P�M�th���(h���!^��]� �E�P�E�   �E�D�h���M�����h�n�E�P�1� h������h�n�E�P�� h���s���h�n�E�P�� �����U���(�H�3ŉE�S�ًM���u3�[�M�3���� ��]� �C V�W��t3�s0�>�;�s'�G���K _�^�B��E�[�M�3��� ��]� �{P u_^���[�M�3��k� ��]� �S�CD9u�C8�K<��C��C,+ɉ�M�{@ u-�sP��P�� �����;�EM_^��[�M�3��� ��]� �M�   �E� W�f�E�E��CE�M��E�   �@ ���    �}��s@�E܋>P�E�M�CM�U�CU��PR�E�P�E�P�E�P�CHP���W����   ��a�}��M�u܃��E�C�+�t�sP�E�V��C�jP�� ��;�uO�E��CE9E�u���v����}� s5Vj�M��5����`����]�#��u�sP�u�������������EM�������}�r�u��
$  ���M�_^��3�[��� ��]� �̃��� ����������U���V��F<�t
���^��]� S�]���u
[3�^��]� W�t#�F ���t�~8;�s�F0��F ʉ8�F0+ω�F ���t*�~0��;�sI��V _�2�ÍN�
�[^��]� ��u3���F0�N�8+9������ s�    ���t�d$ ����+�;�s��u��u_[���^��]� �9P�N@�E��B����N�؋	�M���tWQS��� �M�����u@�F�U��}��^8��F ��F0��F�F<��Ft�     �F,��u��F,�    �h�}���+�F8�F �+ыN��+��F Ӌˉ�F0+�M���F<t�F��F�     �F,�� �F ��F��F+ω�Fˉ�F,+�B��F<t	W�."  ���F0�N<��N _�[�B��E�^��]� ����������U��S�]V��F���t,�F9s%���t�A�;�u�F,� �F^�3����E�[]� �FP��t8���t3�~@ u��PQ�k� �����u�F�ND9t����J���^��[]� ^���[]� ���������U���V�B�0��t@�B;0v9�M���t:N�t�B<u&�B,� �B����t�B^� ���]� 3ɋ�^]� ���^]� ���������U��V��W�F�};�s1�;�w++���;Fu	j���&����N��t*�����F_^]� ;Fu	j��� ����N��t���F_^]� �����������U��V��W�N�};�sF�;�w@+�����*���������;Nu	j���H����N��t3����P�����F_^]� ;Nu	j�������N��tW������F_^]� ����U��V��W�N�};�s=�;�w7+�����*���������;Nu	j����������ȋN��t7j�j P�;Nu	j�������N��tj�j W�A   �A    � �����F_^]� ��������U��j�h��d�    P��SVW�H�3�P�E�d�    �e��ى]�{��+���Q��������ʋu;�v)i��   3WV�EP��������M�d�    Y_^[��]� s��+�P��������E�    �{�EP��+���Q��������ʋ�+�PW�|������E������K+���Q���������+�i��   s�M�d�    Y_^[��]� �M������j j �� ������������U��j�h��d�    P��SVW�H�3�P�E�d�    �e��ى]�s��+;��������������ʋ};�v-����+ǋ��VP�EP���V����M�d�    Y_^[��]� s��+�P���d����E�    �EP���  ��+�Q�s�������E������s��+���������������+�����+ǍƉC�M�d�    Y_^[��]� �M��6���j j �� ������������̋A�8 t�Q,���~H��I��B��Ë�`���������U��SV��W�F�ND9u�}u�~@ u�}�]��������]�}�~P ��   ���]�����tz��ËEu��tPSW�vP��� ����uZ�EP�vP�G� ����uG�V�FD9u�F8�N<��F��F,+ɉ�E�M�H�M_�H�NH^�     �@    �H[]� �E�H_��L^�H�@    �@    �@    []� ���������������U��E�H��L�H�@    �@    �@    ]� U��QS��V�S W���t9C8s�C8�M����   �C�0�u�����   �E��u�K�C8+�u�}����6��u��u�K�}��+�u������t�5H�=L��}�u���
  ���   �C��C8+��;���   |;���   +M��C,�)�C�E��   �C � �E����   �C��C0��C M��C0+ʉ�   ����   ��U��t~�E��u�K�C8+�u�}����1��u�K�u�}��+������t�5H�=L��}�u��|8��r2�C��C8+��;�#|;�w+M�C0�)�C ��u�}���t�5H�=L�E�x_�0^�@    �@    �@    [��]� ���U����ES�]V��E��~P �EW�}�E���   �t�����tw�E�P�vP��� ����ud���tjSW�vP��� ����uK�E�P�vP�R� ����u8�E�ΉFH�T����E�M��H�M�_�H�NH^�     �@    �H[��]�  �E�H_��L^�H�@    �@    �@    [��]�  �������U��E�H��L�H�@    �@    �@    ]�  U��QS�]V�uuW]���W ���t9G8s�G8�L;5Hu;���   �M$��tt�G� �E���tc��|W��rQ�G��G8+��;�B|;�w<+M��G,�)�G�E$tx�G � �E$��tl�G��G0��G M$��G0+ʉ�Q�L�C�L��t7�: t2��|���rߋG��G8+��;��|;�wʋG +�G0�)�G ��؋5H�E_�0^�X�@    �@    �@    [��]�  ���������������U��V��NP��t;�U��u�EEu�B�3��uPRQ�#� ����uj�vP��������^]� 3�^]� ̋�� �����������U��U��t�Ay8 u���E]����]� ����������̋A���t�A,�8 ~�Ë�`������3�3�������������V�q+1���������������^������V��F� ��t;�N,���~�B���F�A��^Å�t�N,���~H��N��B�������P���u�^ËF���t�F,�8 ����^�`V��~P t �j��P���t�vP��� ����y���^�3�^����U���(�H�3ŉE�S��V�C���t.�S,�2�;�s"�F���K^�[�B���M�3��6� ��]Ã{P u^���[�M�3��� ��]ËS�CD9u�C8�K<��C��C,+ɉ�{@ u#�sP�q� �����t�^��[�M�3���� ��]�W�sP�E�   �E�    �E� �;� �������   Pj�M������}��K@�E؋P�E�P�E�P�E�P�E�}�C}�u�Cu��PV�CHP�R��xi��~-��u_�}�rE�}��E�CE�jP�E�jP��� ���u��:�E�9E؋E�uS�}��M�CM�+�Pj �M��u����sP�� ������S�������}�_r�u���  ���M���^3�[��� ��]Ã}��u�Cu�+�u��~���    �D��sPNP�w� �����h����E����V���P���u�^ËF,��N^��B��������������V��F���t�F,� �;�s�^ËW���P�����u_�^ËW���P��_^���̃���������������V�q���u���^�W�y,��;�s�_^��A<u,�A � ��t#;�w9Q8v9A8s�A8�A8+��A_� ^� �_���^��������U���S�]W�W�M�fE�����   �}����   �U�E��U�E�V�c������E��|L��tF;�|;�s���]��t�M�V�A�0�u�^� ��uu��E�M�E+�؋A,)0�A0�(�M���P���t-�MA�E��A��M�U �M����������t���|���j����U�E�^_[��]� �U�E�_[��]� �����U���S�]W�W�M�fE�����   �}����   �U�E��U�E�V��������E��|L��tF;�|;�s���]��t�M�V�A �u�0�n� ��uu��E�M�E+�؋A0)0�A 0�)�u�M���P�R���t'�M�F�E��u�U ���������s���|���i����U�E�^_[��]� �U�E�_[��]� �����k   ��������������������������U��E�� tHt3�]ù̴��J �����]ø   ]������j j j jdjdhZ� j���M  � ����U���VWhp�jjH�j  ������t���Z �O�L��̸���3�����M�@Q�@�С��j �@j��@�M�h��Q��������E��$P�M��Qq �0Wj�K ��PVj j�K ��PhZ� �;u ���M�����r ����E�IP�I�у���_^��]��U��V��N�R�������Y �Et	V�  ����^]� �����jh��������tF� ��@@    �@D    �@H    �@L    �@P    �@T    �@X    �@\    �@`    �3�����������U��M��t�j�P]�����������������A@    �AD    �AH    �AL    �AP    �AT    �AX    �A\    �A`    �����������V�����FX��tP��������FX    �F\    �F`    �FL��tP�������FL    �FP    �FT    �F@��tP�������F@    �FD    �FH    ���^�U��]��  �������U��U�E�M�Z�p�(��"f(��\��\�f(��\��Y��A�\��Y�W��\�f/�rf�E(��8�\A�H�\I(��\�Y�(��\�Y��\�W�f/�r*�\X�\p�\��\��Y��Y��\�f/�r�]� 2�]� U�������*V�qL�IP+�����W�����W҅�~>�O�3��I�����$    �d$ �L0�0�Y1�YD1�ȃ��\��X�Ou��Y(�_^�U��E���]�����U����ESVW�}����^L�@�E���@�E�ˋ��d��\��\d��@�t��<�(��\�f(��\L��]��e��Y��Y��\��Ff/�v_^2�[��]� �}3�����   �EW��;���   ;u��   ;u��   �Ef(ǋ��\ˍ@�\��$�f(��\T�f(��\��Y�f(��\D��Y��\�f/�rX���L�f(��\��\��\��Y�f(��\��Y��\�f/�r#�\\��\$��Y]��Ye��\�f/��"����EF;��6���_^�[��]� �����������U���<SW������*�WP+WL�}���������ڃ��  3ɋú   ����V���Q�:��������ωu��E� �����]��E�3�f/ �v]����   ��rAfo@���%  �yH���@��+Ћ����$    �fn�fp� f����� �@;�|�;�}~���A;�|��s��~k��rRfo@���3�%  �yH���@fnË�fp� f�0�+Ћ�fn�fp� fo�f��f�ȃ���@;�|�;�}��+�H����AH;�|��E���S�����  �u���I�M�����  �u�3�;�NЋ�S�Q;�N��E�    �z��;�NE�PR�M�Q�M̉UЉE���������r  �}� �E�M����MЉUԋ��M��Mȋ��F�M��&  �M��U�;�s/�;�w)+����M�;Fuj�������MȋV��t#�����;Fu	j���}����F��t�Mԉ�F�F�M��U�M�;�s8��u�;֋uw,�M�+����M�;Fuj���8����MȋV��t#�����;Fuj�������M��F��t��F�F�M��U�M�;�s?��u�;֋uw3�M�+����M�;Fuj��������MȋV���*  �����  ;F�  j�������M���   �U�M�;�s8��E�;ЋFw,�M�+����M�;Fuj���o����MȋV��t#�����;Fuj���N����M��F��t��F�F�M��U܉M�;�s8��u�;֋uw,�M�+����M�;Fuj���	����MȋV��t#�����;Fuj��������M��F��t��F�F�MԍU؉M�;�s��u�;֋uw�M������;Fuj�������MԋF��t��F;�}�M���D��G;�|�K���M��UЃ��.����u�V�u�����^_[��]� ���������U��Q�u�E�j P�u�u�u�   ����]� ������������U��j�h��d�    PQSVW�H�3�P�E�d�    �e��E�    �]�u�}��$    ;�tWS�M�B   ���]���}���E������ËM�d�    Y_^[��]�j j �l� ����������������U��M��t�E�~ f��~@f�A�~@f�A]� ���U��V���u����Et	V�Y�������^]� ���������������U���EV�����t	V�(�������^]� ��������������U��j�h��d�    P��SVW�H�3�P�E�d�    �e���3��u�}��t%�����
w���P���������u��u�ܝ �E�    V�s�3���>����E������K+����*��������ʉM���tP�r������M��ƉC�I�ƉC�3�M�d�    Y_^[��]� �u��<�����j j ��� ����������������U��S�YV�q��+ָ���*��������W�}�;�sh+1����*��������򸪪�
+�;�rQ+����*�������������꿪��
+�;�s3�;�_B�^[�E]�����;�_B�^[�E]����_^[]� h���ڜ ���������������U���EZ�����D$�EZ��D$�EZ��$�P]� ��������U����A@�]�U�M�]��U��M�;ADu0f�Yf�Y(f�Qf�Q0�E�f�I f�I8P�I@�
  ��]� �Af/�v�Y�Af/�v�Q�A f/�v�I f/Y(v�Y(f/Q0v�Q0f/I8v�I8�E�P�I@�   ��]� ��������������U��E�I@�@�E��fZ�� �D��EfZ�� �D��EfZ�� ]� ��������������U��E�I@�@�E��� �D��E� �E�D�� ]� ����������U��V��W�N�};�s\�;�wV+�����*���������;Nu	j���x������ȋF��tW�~f� �~Af�@�~Af�@�F_^]� ;Nu	j���5����F��t�~f� �~Gf�@�~Gf�@�F_^]� �������̋A@�AD�AL�AP�AX�A\��������������U���(�E�EV���     �F�F@�u�;FD�L  �FL�NLS�A�F(�N0�\F�\N�V8�\V W�M�f/�v$f/�vf/��E    v�   �I�   �{��Df/�v#f/�vf/��E   v3ۍ{�$�   3��f/��E   v3ۍ{�3��   �F@�ND�E�+ȸ���*��������E�tR�M��E�<��ٍ4��	��$    ����M��E���E���E�P�E��	����M��v�[�uˋu��FX�~XW�ΉG�����O+���������E��t�_[^��]� _[3�^��]� 3�^��]� �%��%��%��%���������U�졠��@���  ]��������������U�졠��@���   ]��������������U�졠��@��  ]���������������+  �����������U�����E��t;�} �u�I�u�   t;�B�P���   �Ѓ�]Ã�B�P���  �Ѓ�]ù   ;�VB�W�xW�R� ������u_^]À} tWj V脴 �������_�F���   ^]�����������U��M��t+�=�� t�y���A�u	�E]�� ����@�M� ]��]����������U��M��t����@�M��@  ]��]á��hﾭދ@��@  ��Y����������U��V�u���t���Q�@� �Ѓ��    ^]�����������U�졠��@���  ]��������������U��E��t�x��u�   ]�3�]������U�졠��@��  ]�������������̡���@��   ��U��E�   ;�VB�W�xW��� ������u_^]À} tWj V�	� �������_�F���   ^]���������������̡���@$�@X�����U�졠��@$�@\]�����������������U���u����u�@$�u�@`Q�Ѓ�]� ��������������̡��V�@��@V�С��V�@$�@D�Ѓ���^�����������U�졠�V�@��@V�С��V�@$�@D�С���u�@$V�@d�Ѓ���^]� ���U�졠�V�@��@V�С��V�@$�@D�С���u�@$V�@�Ѓ���^]� ���U�졠�V�@��@V�С��V�@$�@D�С��V�@$�u�@L�Ѓ���^]� ��̡��V�@$��@HV�С��V�@�@�Ѓ�^�������������U�졠��u�@$Q�@L�Ѓ�]� �����U�졠��@$�@]����������������̡��Q�@$�@�Ѓ����������������U�졠����@$V�@WQ�M�Q�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]� ���U�졠��u�@$Q�@�Ѓ�]� �����U�졠����@$V�@ WQ�M�Q�Ћ���}�IW�I���ы��W�A$�@D�С��W�@$V�@L�С���H$�E�IHP�ы���E�IP�I�у� ��_^��]� ����U�졠����@$V�@$WQ�M�Q�Ћ���}�IW�I���ы��W�A$�@D�С��W�@$V�@L�С���H$�E�IHP�ы���E�IP�I�у� ��_^��]� ����U���,�E�VWP�o������P�I$�E�P�A�Ћ���}�IW�I���ы��W�AV�@�С���M��@Q�@�С���H$�EԋIHP�ы���EԋIP�I�у� ��_^��]� ������̡��Q�@$�@(��Yá��Q�@$�@h��Y�U�졠��u�@$Q�@,�Ѓ�]� �����U�졠��u�@$Q�@0�Ѓ�]� �����U�졠��u�@$Q�@4�Ѓ�]� �����U�졠��u�@$Q�@8�Ѓ�]� �����U�졠��u�@$�u�@PQ�Ѓ�]� ��U�졠��u�@$Q�@T�Ѓ�]� �����U�졠��@$�@l]����������������̡���@$�@p�����U�졠�V�@$��@LV�u�Ѓ���^]� ���������������U�졠�V�@�u�@V�С��V�@$�@D�С��V�@$�u�@L�Ћ���u�I$V�I@�у���^]���U�졠�V�@$�u�@@��V�Ѓ���^]� ���������������U�졠��u�@$Q�@<�Ѓ�]� �����U�졠��u�@$Q�@<�Ѓ����@]� U�졠����@$V�@tWQ�M�Q�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]� ��̡���@$�@x�����U�졠��@(�@]����������������̡���@(�@�����U�졠��@(�@]�����������������U�졠��@(�@]�����������������U�졠��@(�@ ]�����������������U�졠�j�u�@(�u�@��]� ����U���u����u�@(�u�@$��]� ��̡���@(�@(����̡���@(�@,����̡���@(���   �ࡠ��@(�@0�����U�졠��@(�@4]�����������������U�졠��@(�@X]�����������������U�졠��@(�@\]�����������������U�졠��@(�@`]�����������������U�졠��@(�@d]�����������������U�졠��@(�@h]�����������������U�졠��@(�@l]�����������������U�졠��@(�@p]�����������������U�졠��@(�@t]�����������������U�졠��@(�@x]�����������������U�졠��@(���   ]��������������U�졠����@V�@��M�Q�Ѓ��E�P���   ��u3������M��@$Q�u�@�Ѓ��   ����E��IP�I�у���^��]� ������U��Q����U��@(R�@X�Ѕ�u��]� �E3�8M�����   ��]� ���������U������W���E�    �@(�M��@hQ���Ѕ�u_��]� �E���uE����M�@Q�@�С���u�@�M�@Q�С���M�@Q�@�Ѓ��   _��]� �V�ȋ�;���   ;���   h �hx  Q�o���������tg���j �A(�u��@V���Ѕ�u�EP�u������3�^_��]� ���j �H�E�HP�AV�u�ЍEP�u�O������   ^_��]� ���j��@(�ϋ@4��^3�_��]� ����U�졠�V�@(W�}�@pW���Ѕ�t9����΋P(�GP�Bp�Ѕ�t"����΋P(�GP�Bp�Ѕ�t_�   ^]� _3�^]� ���U�졠�V�@(W�}�@tW���Ѕ�t9����΋P(�GP�Bt�Ѕ�t"����΋P(�GP�Bt�Ѕ�t_�   ^]� _3�^]� ���U�졠�S�@(V�@pW�}W���Ѕ���   ����΋P(�GP�Bp�Ѕ���   ����΋P(�GP�Bp�Ѕ�to����_�@(S�@p���Ѕ�tX����΋P(�CP�Bp�Ѕ�tA����΋P(�CP�Bp�Ѕ�t*�GP��������t�G$P��������t_^�   []� _^3�[]� �����U�졠�S�@(V�@tW�}W���Ѕ���   ����΋P(�GP�Bt�Ѕ���   ����΋P(�GP�Bt�Ѕ�to����_�@(S�@t���Ѕ�tX����΋P(�CP�Bt�Ѕ�tA����΋P(�CP�Bt�Ѕ�t*�G0P���-�����t�GHP��������t_^�   []� _^3�[]� �����U�졠��@(�@8]�����������������U�졠��@(�@<]�����������������U�졠��@(�@@]�����������������U�졠��@(�@D]�����������������U�졠��@(�@H]�����������������U�졠��@(�@L]�����������������U�졠��E�@(Q�@P�$��]� �U�졠��E�@(���@T�$��]� ���������������U�졠��u�@(�u�@|��]� ������U�졠��u�@(�u���   ��]� ���U�졠��� �@$V�@W�u���M�Q�Ћ�����I�E��IP�ы���A�M��@QV�С���M��@Q�@�Ѓ��E�P���L   ������I�E��IP�у���_^��]� �����������U�졠��} �P(�����E�B8]����U�졠�S�@V�@dW�ًMj �Ѝx�Ǚ�ȋ�;�u|;�uxh �h�  Q�C���������t_����M�Bj �@hWV�С��W�@(�ˋ@H�Ѕ�t���W�@(V�@ ���Ѕ�t�   �3��EP�u�'�������_^[]� ���j��@(�ˋ@4��_^3�[]� �U�졠�V�@(W�}�@P�Q���$�Ѕ�tG����G�@(Q�@P���$�Ѕ�t)����G�@(Q�@P���$�Ѕ�t_�   ^]� _3�^]� ������������U�졠�V�@(W�}�@T������$�Ѕ�tK����G�@(���@T���$�Ѕ�t+����G�@(���@T���$�Ѕ�t_�   ^]� _3�^]� ������U�졠�V�@(W�}�@P�Q���$�Ѕ��  ����G�@(Q�@P���$�Ѕ���   ����G�@(Q�@P���$�Ѕ���   ����G�@(Q�@P���$�Ѕ���   ����G�@(Q�@P���$�Ѕ���   ����G�@(Q�@P���$�Ѕ�tt����G�@(Q�@P���$�Ѕ�tV����G�@(Q�@P���$�Ѕ�t8����G �@(Q�@P���$�Ѕ�t�G$P���������t_�   ^]� _3�^]� �����U�졠�V�@(W�}�@T������$�Ѕ���   ����G�@(���@T���$�Ѕ���   ����G�@(���@T���$�Ѕ���   ����G�@(���@T���$�Ѕ�ti����G �@(���@T���$�Ѕ�tI����G(�@(���@T���$�Ѕ�t)�G0P���R�����t�GHP���C�����t_�   ^]� _3�^]� �����������̡���@(� ������U�졠�V�@(�u�@�6�Ѓ��    ^]���������������U�졠��@(���   ]��������������U�졠��@(�@]����������������̡���@(�@�����U�졠�V�@(�u�@�6�Ѓ��    ^]���������������U�졠��u�@,�u�@Q�Ѓ�]� �̡���@,�@����̡���@,�@����̡���@,�@����̡���@,�@ ����̡���@,�@(����̡���@,�@$�����U�졠��@,�@]�����������������U�졠����@,V�@W�U�R�Ћ���}�IW�I���ы��W�A$�@D�С��W�@$V�@L�С���H$�E�IHP�ы���E�IP�I�у���_^��]� ����̡��j �@,j � �Ѓ��������������U�졠�V�@,�u�@�6�Ѓ��    ^]��������������̡���@,�@4����̡���@,�@8�����U�졠����@,V�@<W�U�R�Ћ���}�IW�I���ы��W�A$�@D�С��W�@$V�@L�С���H$�E�IHP�ы���E�IP�I�у���_^��]� �����U�졠����@,V�@@W�u�U�R�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]� ̡���@,�@,�����U�졠�V�@,�u�@0�6�Ѓ��    ^]���������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@�@]�����������������U�졠��@�@]�����������������U�졠��@�@]�����������������U�졠��@�@]�����������������U�졠��@�@]�����������������U�졠��@�@]�����������������U�졠��u�@�u�@\��]� ������U�졠��u�@�u��  ��]� ���U�졠��E�@���@ �$��]� ���������������U�졠��E�@Q�@$�$��]� �U�졠��E�@���@(�$��]� ���������������U�졠��@�@,]�����������������U�졠��@�@0]�����������������U�졠��@�@4]�����������������U�졠��@�@8]�����������������U�졠��@�@<]�����������������U�졠��@�@@]�����������������U�졠��@�@D]�����������������U�졠��@�@H]�����������������U�졠��@�@L]�����������������U�졠��@�@P]�����������������U�졠��@���   ]��������������U�졠��u�@Q��  �Ѓ�]� ��U�졠��@�@T]�����������������U�졠��@�@X]�����������������U��U��u3�]� ���R�@ Q�@(�Ѓ��   ]� �����U�졠��@���   ]��������������U�졠��@��  ]��������������U�졠��@�@`]�����������������U�졠��@�@d]�����������������U�졠��@�@h]�����������������U�졠��@�@l]�����������������U�졠��@�@p]�����������������U�졠��@�@t]�����������������U�졠��@���   ]��������������U�졠��@��  ]��������������U�졠��@�@x]�����������������U�졠��@�@|]�����������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��u�@Q��  �Ѓ�]� ��U�졠��@���   ]��������������U�졠��@���   ]��������������U��U��t���R�@ Q�@$�Ѓ���t	�   ]� 3�]� �U�졠�Q�@ �u�@L�u�Ѓ�]� ��U�졠��@���   ]��������������U�졠��@��  ]�������������̡���@���   ��U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]�������������̡���@���   ��U�졠��@���   ]�������������̡���@���   �ࡠ��@���   �ࡠ��@��   �ࡠ��@���   ��U�졠��@��  ]�������������̡���@���   �ࡠ��@���   ��U�졠�V�@�u���   V�Ѓ��    ^]�������������U�졠��@� ]�ࡠ��@�@�����U�졠��@���   ]��������������U�졠��@��   ]��������������U�졠��@�@]�����������������U�졠��@�@]�����������������U�졠��@�@]�����������������U�졠��@�@]�����������������U�졠��@�@]�����������������U�졠��@���  ]��������������U�졠��@�@]�����������������U����E�V�uP����������M�@$Q�@�Ѓ���t]����M�@j�@Q�Ѓ���u�E�P��������t3���j�@V�@�Ѓ���u���V�@�@�Ѓ���t�   �3�����H$�E�IHP�ы���E�IP�I�у���^��]��������U�졠��@�@ ]�����������������U�졠��@�@(]�����������������U�졠��@��  ]��������������U�졠��@��   ]��������������U�졠��@��  ]��������������U�졠��@��  ]��������������U�졠����@V�@$�M�WQ�Ћ���}�IW�I���ы��W�A$�@D�С��W�@$V�@L�С���H$�E�IHP�ы���E�IP�I�у���_^��]��������U�졠����@V���  �M�WQ�Ћ���}�IW�I���ы��W�A$�@D�С��W�@$V�@L�С���H$�E�IHP�ы���E�IP�I�у���_^��]�����U��j�u�  �E��]������������U���<��SVW�E�    ��t�E�P�   �h������-����M��@Q�@�   �С���M��@$Q�@D�Ѓ��}ࡠ��u�@V�@�С��V�@$�@D�С��V�@$W�@L�Ѓ���t(����M��@$Q�@H����С���M��@Q�@�Ѓ���t&����H$�EċIHP�ы���EċIP�I�у�_��^[��]������U�졠����@V���  W�u�M�Q�Ћ���}�IW�I���ы��W�A$�@D�С��W�@$V�@L�С���H$�E�IHP�ы���E�IP�I�у� ��_^��]��U�졠��@��D  ]��������������U�졠��@��H  ]��������������U�졠��@��L  ]��������������U�졠����@V���  W�u�M��uQ�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]��������������U�졠��@���  ]��������������U�졠��@���  ]�������������̡��V�@j �@j����Ћ�^���������U�졠�V�@j �u�@���Ћ�^]� �U�졠�V�@�u�@j����Ћ�^]� ̡���@�@�����U�졠�V�@j ���   ��Mj V�Ћ�^]� �����������U�졠��u�@Q�@�Ѓ�]� �����U�졠��u�@Q�@�Ѓ����@]� U�졠�h#  �u�@�u�@l��]� �U�졠�hF  �u�@�u�@l��]� �U�졠��u�@�@t�Ћ��P���   �@X�Ѓ�]� ����U�졠��u�@�@t�Ћ���u�Ћ��   R�@`�Ѓ�]� ���������������U�졠��u�@���   �Ћȅ�u]� ���Q���   �@�Ѓ�]� ��������U�졠��@���   ]���������������l��A    �A    �A    �����V��~ �l�u����v�@4� �Ѓ��F    �F    ^���������������̸   ����������̸   �����������3�� ������������ �������������U�졠�V�@4��@$h�  �v���u����u�@4�u�@�u�v�Ѓ�2�^]� ���������������U���u��u�u�u�P]� ��������3�� ����������̸   � ��������� �������������U��Q���S�@V�@ W�}�ًω]�3���=INIb�  ��   =SACbmt)=$'  t
=MicM�f  �W���P$�   _��^[��]� ��MQ�M�Q�ˉu��u�P��t�u����u��@4�s�@�Ѓ��   _��^[��]� =ARDb�  ���j �@j���   ���Ћء��j �@j���   ���ЋM�����j �@j���   �ЋM�𡠴j �@j���   ���u�M�P�VWS�R�   _��^[��]� ����P�   _��^[��]� =NIVb_tF=NPIbt.=ISIbuV�3���  P���r  P���V�   _��^[��]� �W���P_^[��]� ����P�   _��^[��]� =cnyst_��^[��]� ���j �@hIicM���   ���ЋWP���R _^[��]� �������U���,V��~ t~����v�@4�@�Ѓ} t���P�F�I0�p�Al�Ѓ�^��]� ���M�hARDb�E��E�    �����NP�E�P�E�P�  ����M苀�   Q� �Ѓ��M�����^��]� ������������U�졠��u�@4�q�@l�Ѓ��   ]� �������������̡���q�@4�@�Ѓ�������������̡���q�@4�@�Ѓ�������������̡���q�@4�@�Ѓ�������������̡���q�@4�@|�Ѓ�������������̡���q�@4���   �Ѓ�����������U�졠��u�@4�q�@(�Ѓ�]� ���U���u����u�@4�u�@,�q�Ѓ�]� �������������U���u����u�@4�q�@0�Ѓ�]� ����q�@4�@4��Y���������������U�졠��u�@4�q���   �Ѓ�]� U�졠��u�@4�q�@ �Ѓ�]� ���U�졠��u�@4�q�@$�Ѓ�]� ���U�졠�V���   �u�@WV���Ѓ������V���   u �@@�Ћ��P�I4�w�A �Ѓ�_^]� �@�Ѓ���u,���V���   �@8�Ћ��P�I4�w�A$�Ѓ�_^]� hh�h�  hx�h  @��  ���=�� t
�=�� t�_^]� ���U���u����u�@4�q�@D�Ѓ�]� U���u����u�@4�q�@H�Ѓ�]� U���u����u�@4�q�@L�Ѓ�]� U���u����u�@4�q�@P�Ѓ�]� U�졠�S���   V�@W�}W���Ѓ���������   �@��   �uV�Ѓ������V���   u6�@@�Ћ��W���   ���I@�ы��V�I4P�s�AP�Ѓ�_^[]� �@�Ѓ���uB���V���   �@8�Ћ��W���   ���I@�ы��V�I4P�s�AH�Ѓ�_^[]� hh�h   ��   W�Ѓ�����   ����u���   V�@�Ѓ������V���   u6�@@�Ћ��W���   ���I8�ы��V�I4P�s�AL�Ѓ�_^[]� �@�Ѓ���uB���V���   �@8�Ћ��W���   ���I8�ы��V�I4P�s�AD�Ѓ�_^[]� hh�h)  �
hh�h-  hx�h  @��  ���=�� t
�=�� t�_^[]� ��������������U���u����u�@0�u���   �u�q�Ѓ�]� �������U�졠��u�@0�q���   �Ѓ�]� U���E������@0�$�u���   �u�q�Ѓ�]� U���u����u�@4�u�@�u�q�Ѓ�]� ����������U���u����u�@4�u�@�u�q�Ѓ�]� ����������U���u,����u(�@4�u$�@T�u �u�u�u�u�u�u�q�Ѓ�,]�( ��������U���u����u�@4�u��  �u�q�Ѓ�]� �������U���u$�E�u ����u�@4�u��  ���D$�E�$�q�Ѓ�$]�  ���������������U�졠�h�����@4h�����@Th�����u�uh����h����h����h�����u�q�Ѓ�,]� ����������U�졠��u�@4�q�@8�Ѓ�]� ���U�졠��u�@4�q�@<�Ѓ�]� ���U���u����u�@4�q���   �Ѓ�]� ������������̡���q�@4�@@�Ѓ�������������̡���q�@4��  �Ѓ�����������U�졠��E�@4����  �$�q�Ѓ�]� ������U���u����u�@4�u�@X�u�q�Ѓ�]� ���������̡���q�@4�@`��Y��������������̡���q�@4�@d�Ѓ��������������U���u����u�@4�u��   �u�q�Ѓ�]� �������U���u����u�@4�u�@\�u�u�u�q�Ѓ�]� ���̋I��u��á��Q�@4��   �Ѓ���U���u����u�@4�q��  �Ѓ�]� �������������U���u����u�@4�q�@h�Ѓ�]� U���u����u�@4�q��  �Ѓ�]� �������������U���u����u�@4�q�@p�Ѓ�]� U���V��hYALf�M���������P�R4�v�Bl�Ѓ��M�����^��]���������U��QVW�}�M���t����M�@j ���   j�Љ�u��t����M�@j ���   j�Љ����M��@4V�@pW�q�Ѓ�_^��]� �������U���u����u�I�@0�u���   �q�Ѓ�]� �������U���u����u�@4�u�@x�u�q�Ѓ�]� ����������U�졠��u�@4�q�@t�Ѓ�]� ���U���u����u�@4�u���   �u�u�q�Ѓ�]� ����U���u����u�@4�u���   �u�u�q�Ѓ�]� ����U������SW�E�    �E�    �@�ًM���   �{j j�ЋM�E����j �@j���   �ЉE�����M��@0Q�@`�M�Q�w�С���s�@4�@�Ћ��j �I0�U�R�U�R�U�R�U�RP�C�p�Ah�Ѓ�,�} _[t(�} t(�M�U�;�~<�E��;�}3�M��U�;�~)�E���} u�M�U�;�~�E��;�}�   ��]� 3���]� ���U���u�E������@4�D$�E���   �$�u�q�Ѓ�]� �����U���u����u�@4�u���   �q�Ѓ�]� ���������̡���q�@4���   �Ѓ����������̡���q�@4��  �Ѓ�����������V��V������h���@0� �Ѓ��F�F    ��^�����V��N�����t���Q�@0�@�Ѓ��F    ^������̸   ����������̸   ����������̸   � ��������3�� �����������3���������������� �����������������������������U�졠�V�@W�}�@ �����=NIVb��   ��   =TCAbwtM=$'  t3=MicM��   ���j �@hIicM���   ���ЋWP���R_^]� �W���P_�   ^]� ���j �@hdiem���   ���ЋWP���R_^]� =INIbu�~ u�����F   �P_^]� �~ t�����P_^]� =atni@t1=ckhct=ytsdu;����P_�F    3�^]� ����P_^]� �5  _3�^]� =cnys����_3�^]� ����������U��V��N��u3�^]� ���j �@0j ���   j j j �u j �ujQ���u����u�@0�u���   �uj �u�v�Ѓ�D^]� ����������̋I��u3�á��Q�@0�@�Ѓ�����̋I��u3�� ���Q�@0�@�Ѓ�� U���V�q��u�E�p�    ^��]� �E�H����Q�u�@0R���   �M�VQ�Ћuj �    �F    ���P���   V�I�ы���E����   P�	�у�$��^��]� ��������U�졠��u�@0�q���   �Ѓ�]� ����q�@0���   �Ѓ����������̡��j �@0j ���   j j j j j j j4�q�Ѓ�(�������̡��j �@0j ���   j j j j j j j;�q�Ѓ�(��������U�졠��u�@0�q�@�Ѓ�]� ���U��I��t'���j �@0j ���   j j j j �uj jQ�Ѓ�(]� �����������U���u����u�@4�u�@,�q�Ѓ�]� �������������U���u����u�@4�q�@0�Ѓ�]� ����q�@4�@4��Y���������������U��V�q��u3�^]� �E�H����Q�u�@0R�@V�Ѓ�^]� �����������U��V�q��u3�^]� �E�H����Q�@0R���   V�Ѓ�^]� �����������U��E3�h�����h   ���Pj BRj �u�u�   ]� ���U���$VW��htniv�M��I�������u�@hulav�@4�M��С��hgnlf�@htmrf�@4�M��С���u�@hinim�@4�M��С���u�@hixam�@4�M��С���u�@hpets�@4�M��С���u�@hsirt�@4�M��ЋM �u$��   �u�����t,���Q�@h2nim�@4�M��С��V�@h2xam�@4�M��ЍE�P�u�E�P���S������P���   �@8�Ћ�������   �E��	P�у��M��p���_��^��]�  ������U���$V��htlfv�M��
�������E�@���@,�$hulav�M��С���u,�@htmrf�@4�M��С���E�@���@,�$hinim�M��С���E�@���@,�$hixam�M��С���E$�@���@,�$hpets�M��С���uD�@hsirt�@4�M����U0W�f.џ��Dz�E8f.����D{?������@�$�@,h2nim�M��С���E8�@���@,�$h2xam�M��С���u@�@hdauq�@4�M��ЍE�P�u�E�P���������P���   �@8�Ћ�������   �E��	P�у��M��������^��]�@ ������������U���u,W�j ���D$�$�E$htemf�� �D$�E�D$�E�D$�E�$�u����]�( ��������U���Mf.P�����%�����D{�Y��^��Uf.H����D{�Y��^��u,W�j ���D$�$�E$�Y�hrgdf�� �^��D$�E�L$�T$�$�u�h���]�( ����U���u,���W�j ���D$�$�E$�^�htcpf�� �D$�E�^��D$�E�^��D$�E�$�u�����]�( ����U���0�E�M���u����@���   �Ѕ�u��]� SVW����X  htlfv�MЋ�������u�����yfn���Ƀ��Y��E��E��$�^� �]��F�$�P� �E��]��^E�G,�$hulav�M��С��hmrff�@htmrf�@4�M��Ћu�����xfn���Ƀ��Y��E��E��$�� �]��F�$�ۈ �E��]��^E�G,�$hinim�M��Ћu�����xfn���Ƀ��Y��E��E��$莈 �]��F�$耈 �]��E��^E�G,�$hixam�M��С������@���@,�$hpets�M��С��j �@hdauq�@4�M��С��S�@hspff�@4�M��С���u �@hsirt�@4�M��ЋM��E�P�u�E�P�������P���   �@8�Ћ�������   �E�	P�у��M��1���_��^[��]� ������U���$V��hCITb�M����������u�@hCITb�@8�M��С���u�@hsirt�@4�M��С���u�@hulav�@4�M��ЍE�P�u�E�P���`������P���   �@8�Ћ�������   �E��	P�у��M��}�����^��]� ����U��V�q��u3�^]� �E�E�H����Q�u �@0���@(�D$�E�$�uRV�Ѓ�$^]� U����E�Vj �u��MP�6���P�u�������������I�E��IP�у���^��]� �����������U��V�q��u3�^]� �E�H����Q�@0�M�@,QRV�ЋM3҃�9U^�]� �������������U��V�q��u3�^]� �E�H����Q�u�@0R�@,V�Ѓ�^]� �����������U��V�q��u3�^]� �E�H����Q�u�@0R�@0V�Ѓ�^]� �����������U��VW���O����   �E�P�0���R�u�@0V�@0Q�Ѓ���tf� t`�E�H����Q�p0�E��P�F0R�w�Ѓ���t8���t1�E�H����Q�p0�E��P�F0RW�Ѓ���t_�   ^]� _3�^]� ��������������U��QV�q��u	3�^��]� �E�E�    �H����Q�@0�M��@8QRV�Ћ�����tC�U���t<����u�AR�@�ЋM�����t ���Q�@�@�ЋE��E�EP��������^��]� ���U��V�q��u3�^]� �E�H����Q�u�@0�u�@<RV�Ѓ�^]� ��������U��E��V���u����@���   �Ѕ�u^��]� W����R  �v����t!�E�H����Q�@0�M��@0QRV�Ѓ���fn�������Y���M��D$�E��Y���$�p  �~ �M_f��~@��f�A^��]� �U�졠����@V�@��M�Q�Ѓ��E�P�u���U�������t�M�E�P�#�������E��IP�I�у���^��]� �����U��V�q��u3�^]� �E�H����Q�@0j ���   j j j j j Rj1V�Ѓ�(^]� �������������U�졠�V�@j �u���   ��M��h���h   �j j jj P�u���E���^]� U�졠�V�@j �u���   ��M���u$���u j �u�u�uP�u����^]�  �U������V�@�����   W��$�u��M���]��E8j �u@�΃��D$�E0�$�u,�E$�� �D$�E�D$�E�D$�E��$�u����^��]�< ����U������V�@�����   W��$�u��M���]�j j ��W��D$�$�E$htemf�� ���D$�E�D$�E�D$�E��$�u�1���^��]�$ ����������U������V�@�����   W��$�u��M���]��Uf.P�����%�����D{�Y��^��Mf.H����D{�Y��^�j j ��W��D$�$�E$�Y�hrgdf�� ���^��D$�E��T$�L$�$�u�]���^��]�$ ������U������V�@�����   W��$�u��M���]����j W�j �����D$�$�E$�^�htcpf�� �D$�E�^��D$�E�^��D$�E��$�u����^��]�$ ������U���0���V��W��E�����M�Q�u�E��@�MЋ��   Q�M���~ j �u f�E��u�~@�u�E�P�u���uf�E��U���^��]� ��������������U�졠���0�@V�@W���M�Q�С�����@�M����   Q�u�M�Q�M�Ћ�����I�E��IP�ы���A�M��@QV�С���MЋ@Q�@�Ѓ��E��u��j P�u�����������I�E��IP�ы���A�M��@Q�Ѓ���_^��]� ���U���dV��M��o�������M�RP�u�E�P���   ��P�M�������M��2���j j �E�P�M�貳��P�u���W���������I�E��IP�у��M�������M�������^��]� �������U���P�U���V�uW���E����t+������@W����   �$R�����]��E��E����W��M�Q�u�E��E��E��@�M����   Q�����~ �wf�E��~@f�E��~@f�E؅�u
_3�^��]� �E�E�H����Q�u �@0���@(�D$�E��$�M�QRV�Ѓ�$_^��]� ����U��V�q3���t)�E�H����Q�@0�M�@,QRV�Ћ�3���9E�����P�Q�u�M�R0�ҋ�^]� ��������������U��V�q��t!�E�H����Q�@0�M�@,QRV�Ѓ�������u�A�u�M�@4�Ћ�^]� ������U���V�q��t!�E�H����Q�@0�M��@0QRV�Ѓ�������E��A�M�@,���$�u�Ћ�^��]� �������U���V�E�P�uW��u�E�����E�����������Q�M�R@�E�P�u�ҋ�^��]� ��U���V��W�~W��E��E��E�����   �E�H����Q�@0�M�@0QRW�Ѓ���tx�~��tq�E�H����Q�@0�M��@0QRW�Ѓ���tN�v��tG�E�H����Q�@0�M��@0QRV�Ѓ���t$����M�@Q�u�M�@H��_�   ^��]� _3�^��]� ����U�졠����@V�@��M�Q�Ѓ��E�P�u������������Q�M�R8�E�P�u�ҡ���M��@Q�@�Ѓ���^��]� ��������������U���,V��M��O�������M��@Q�@�Ѓ��E�P�u���-�������u����M��@Q�@�Ѓ�� �E�P�M���������M��@Q�@�Ѓ�����M�P�EԋR<P�u�ҍM��®����^��]� ���������U��� V�qW��E��E��E���t%�E�H����Q�@0�M��@<Q�M�QRV�Ѓ����U���t����A�M��@HQ�MR�ЋU���t����E��@�M�@,���$R�Ћ�^��]� ��������������U��E3҃8V�p�¸   h���h   ���E�3�����Rj @Pj V�u����^]� ��������������U��U�u 3��:�u��P�u�u�u�r�u�W���]� ���U��U�E43��:��P�u<���D$�E,�$�u(�E �� �D$�E�D$�E�D$�B�$�u�-���]�8 ���������U��E3҃8�H��W�Rj ���D$�$�E htemf�� �D$�E�D$�E�D$�$�u�����]�  ���������������U��E�U�h����%��3҃8��f.P����D{�Y��^��Mf.H����D{�Y��^�Rj ��W��D$�$�E �Y�hrgdf�� �^��D$�T$�L$�,$�u����]�  �����������U��E���3҃8W����PRj ���D$�$�E �^�htcpf�� �D$�E�^��D$�E�^��D$�$�u����]�  �����������U��U3��:��P�u�B�u�uP�u�u�i���]� �����U��E�u3҃8��RP�u�r���]� ��������������U���$V��hgnrs�M��*����E�E�����E�   �@�M����   Qj�M��С���M����   Q� �ЋE�E�������E�   �@�M����   Qj�M��С���M����   Q� �Ѓ��E�P�u�E�P���������P���   �@8�Ћ�������   �E��	P�у��M�������^��]� ����U��W�y��u3�_]� �E�E�H����V�p0�EQ�u �����D$�E�$P�F(RW�Ѓ�$^_]� ���������̡��j �@0j ���   j j j j j j j �q�Ѓ�(�������̋I��u��á��Q�@4��   �Ѓ���U��I��u3�]� ����u�@4�u��  Q�Ѓ�]� ��U��I��u3�]� ����u�@4�u�@hQ�Ѓ�]� �����U��I��u3�]� ����u�@4�u�@pQ�Ѓ�]� �����U��I��u3�]� ����u�@4�u��  Q�Ѓ�]� ��U���u����u�@0�u���   �u�q�Ѓ�]� �������U�졠��P0�E�pj j j �u�uj �0���   j=�q�Ѓ�(]� �����������U�졠��P0�E�p�uj j j��uj �0���   j=�q�Ѓ�(]� �����������U��E�u���̴EС���2�@0�u�@@�q�Ѓ�]� �U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   �u�ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   �u�ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u���   �u�u�ujQ�ЋE���(��]� ���������������U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u���   �uj �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u���   �uj �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u���   �uj �uj*Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   j �ujQ�ЋE���(��]� �U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   j �ujQ�ЋE���(��]� �U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   j �uj	Q�ЋE���(��]� �U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   j �uj
Q�ЋE���(��]� �U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u���   �uj �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u���   �uj �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   �u�uj'Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   �u�uj,Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u���   �uj �uj:Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j j �u�E�    �u�@0j ���   j j)Q�ЋE���(��]� ���U��Q�I��u3���]� ����U�Rj j �u�E�    �@0j �u���   j j j)Q�ЋE���(��]� ���U��I��u3�]� ���j �@0j ���   j �u�u�uj �ujQ�Ѓ�(]� ��U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u���   �uj �ujQ�ЋE���(��]� U��Q�I��u3���]� ����U�Rj �u�E�    �u�@0�u���   �uj �uj>Q�ЋE���(��]� U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   j �ujQ�ЋE���(��]� �U�졠�j �@0j ���   j �u�u�uj �uj.�q�Ѓ�(]� �������������U��V�q��u3�^]� �E�H����Q�@0j ���   j j j �u�uRjV�Ѓ�(^]� �����������U��V�q��u3�^]� �E�H����Q�@0j ���   j j j j j RjV�Ѓ�(^]� �������������U��V�q��u3�^]� �E�H����Q�u�@0R�@\V�Ѓ�^]� �����������U���SVW�u�ٍM��
 �EP�E�P�M���
 ��tj�}�I �M��tI���Q���   �@H�ЋS������tN�w���j �A0j ���   j j �u�V�7jR�Ѓ�(��t"�EP�E�P�M��
 ��u�_^�   [��]� _^3�[��]� ���U��Q�I��u3���]� ����U�Rj j �u�E�    �u�@0�u���   j �ujQ�ЋE���(��]� �U�졠�V�@4W�}� �w���ЋE�G    �w�H����Q�u�@0W���   R�v�Ѓ�3Ʌ����G_^��]� �������U��I��u3�]� ���j �@0j ���   j �u�u�uj �uj/Q�Ѓ�(]� ��U��U��u3�]� �r�B    ����u�@0�q���   �Ѓ�]� ���������U��I��u3�]� ���j �@0j ���   j j j �uj j jQ�Ѓ�(]� ����̡��j �@0j ���   j j j j j j j6�q�Ѓ�(��������U��I��u3�]� �u����u�@0�u�@DQ�Ѓ�]� ��U��I��u3�]�  �u$����u �@0�u���   �u�u�u�u�uQ�Ѓ�$]�  �I��u3�á��Q�@0�@X�Ѓ������U��I��u3�]� ����u�@0�u�@LQ�Ѓ�]� �����U��Q��u3�]� ����H0�E   �P�APR�Ѓ�]� ��U��I��u3�]� ����u�@0Q�@P�Ѓ�]� ��������U��I��u3�]� �u����u�@0�u�@T�uQ�Ѓ�]� ���������������U���VW���M��~����E�M�P�0���R�@0Q���   j j j j j Vj8�w�Ћ���(��t�M�E�P�����M�����_��^��]� ����������U��EV�P�0���R�u�@0j ���   j j j j Vj9�q�Ѓ�(^]� ��������U��EV�P�0���R�u�@0�u�@h�u�uV�q�Ѓ�^]� ��������������U��QVW�}�M���t����M�@j ���   j�Љ�u��t����M�@j ���   j�Љ����M��@0V�@`W�q�Ѓ�_^��]� �������U���u����u�@0�u���   �q�Ѓ�]� ����������U��U����@0��t*���   R�q�Ћ���u�ЋA0R���   �Ѓ�]� �u�@|�q�Ѓ�]� ��U���u����u�@0�u�@p�u�u�q�Ѓ�]� �������U���u����u�@0�u�@d�u�u�q�Ѓ�]� �������U�졠�j �@0j �u���   �u�u�uj �uj3�q�Ѓ�(]� ������������U��Ej ����j �@0j ���   j j j j Rj�q�Ѓ�(]� �������������U��Ej ����j �@0j ���   j j jj Rj�q�Ѓ�(]� �������������U��Ej ����j �@0j ���   j j j j Rj�q�Ѓ�(]� �������������U��EV�P�0���R�@0j ���   j j j j j Vj"�q�Ѓ�(^]� ���������U��EV�P�0���R�@0j ���   j j j j j Vj5�q�Ѓ�(^]� ���������U��EV�P�0���R�@0j ���   j j j �uj Vj<�q�Ѓ�(^]� ��������U�졠�V�@0j ���   j j j j �u��j �uj�v�С���u�@0�v�@t�Ѓ�0^]� �������̡��j �@0j ���   j j j j j j j�q�Ѓ�(��������U�졠�j �@0j ���   j j j j �uj j�q�Ѓ�(]� ���j �@0j ���   j j j j j j j�q�Ѓ�(��������U�졠�j �@0j ���   j j j j j �uj�q�Ѓ�(]� U�졠�j �@0j ���   j j j j �u�uj&�q�Ѓ�(]� ��������������̡��j �@0j ���   j j j j j j j(�q�Ѓ�(�������̡��j �@0j ���   j j j j j j j#�q�Ѓ�(��������U�졠�j �@0j ���   j j �u�uj �uj+�q�Ѓ�(]� �������������̡��j �@0j ���   j j j j j j j0�q�Ѓ�(��������U�졠��u�@0�q���   �Ѓ�]� U���V�u ��M��|�������u�@h8kds�@4�M��С���M Q�M�Qj �u�E     �u�@0�u���   �u�uj2�v�Ћu ��(�M��A�����^��]� �������̡���q�@0���   �Ѓ�����������U��I��u3�]� ���j �@0j ���   j j j j j �uj-Q�Ѓ�(]� �����U������W�@j ���   ���Mj�ЋM�E����j �@j���   �ЉE�����M��@0Q�@`�M�Q�w�С���U��H0�E�pR�U�R�U�R�U�R�0�Ah�w�Ѓ�(�} _t(�} t(�M��U�;�~<�E��;�}3�M��U�;�~)�E���} u�M��U�;�~�E��;�}�   ��]� 3���]� �����U��SV�uW��u�q����]�@j ���   hdiuM���Ћ���tI;>u	_^3�[]� ���j �@hIicM���   ����;�u���j �@h1icM���   ���Шu��>_^�   []� ���������U�졠���(�@V�u�@Thfnic���ЋЅ�t���j
�A�ʋ��   �Ѕ���   ���hfnic�@�M؋@PQ����P�M��޸���M�������u�E�P��������M���������΋@�@ �Ѓ��t����΋@�@ �Ѕ�u���hfnic�@�΋@$�С���u�@j
�@8����^��]������������̡���q�@0���   �Ѓ�����������U���$V��hmnrs�M��
�������u�@j�@4�M��ЍE�P�u�E�P����������P���   �@8�Ћ�������   �E��	P�у��M�������^��]� �������U���$�} V��SSSS�DSSSE�P�M��}�������M܋@�@ �Ћ��j�QP�B4�M��ЍE�P�u�E�P���7������P���   �@8�Ћ�������   �E��	P�у��M��T�����^��]� �����������V��V������h���@0� �Ѓ��F�F    ����F   �F    ��^�V��N�����t���Q�@0�@�Ѓ��F    ^�������U��V��N�F    ��tg���j �@0j ���   j j j j j j jQ�С���u�H0�u3�9E�u���uj ��
P�v���   �Ѓ�D��t�~ t
�   ^]� 3�^]� ��������������U��E�A�I��u3�]� ���Q�@0�@�Ѓ�]� �����U�졠�S�@�]�@ V�����=ckhc��   t|=cksatb=TCAb��   ���W�@j ���   hdiem���Ћ��SW���F   �R�~ ��t��t��u3�������P�J���_^��[]� �~ ti����P^[]� �~ tV���j �@0j ���   j j j j j j j �v�Ѓ�(��t*�F    ^�   []� =atnit�u��S�����^[]� ^3�[]� ����������U��Q�y �M���   S�]V�uW�}��wp�$���9u��   �^9u��   �S9u��   �H9u��   �=�E;�~6;���   �,�E;�|%;�~}��E;�|;�|p��E;�~;�~c�9uu\���j �@0j ���   j j j j j �uj�q��fn������(j���D$fn�����$S�oJ  �E����@    _^[��]� ������������� �-�����U��W��� �6  V�u����   �$���Ef/E�  �   �Ef/E��   �   �Mf/M��   �   �Mf/M��   �|�Uf/Uvp�E f/���   �_�Uf/UrS�E f/���   �B�Uf/Ur6�E f/�w�)�Uf/Uv�E f/�sf��Ef.E���DzT���j �@0j ���   j j j j j �uj�w���E ��(�u(���D$�E�$V��H  ���G    ^_]�$ ������#�5�R�o�����U���E j���D$�E�D$�E�$�u�u�]���]�  ���������U���E j���D$�E�D$�E�$�u�u����]�  ���������U���E j���D$�E�D$�E�$�u�u�����]�  ���������V��V������h���@0� �Ѓ��F�F    ����F   ��^��������V��N�����t���Q�@0�@�Ѓ��F    ^�������U�졠�V�@��M�@ ��=cksat]=ckhct�u���u�����^]� j j j j j j �F   ���j �@0j ���   j �v�Ѓ�(��t#�F    �   ^]� �~ t����P^]� 3�^]� �������������U��V��V������h���@0� �ЋM�F�E�F    �F   ���F������@j ���   hmyal�ЉF��t��t�F    ����M�@j
���   hhfed�ЉF��^]� U�졠�V�@��M�@ ��=ytsdt�u���u����^]� ����v�@0���   �Ћ�����P�   ^]� ����������3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U���V�u�E�    �V�E�    �    �B    ��������j ���   �E��IPR�ы���E����   P�	�у���^��]� ����������̋A��uË ���������������������U��V���PD��t�E9Ft
�F����PH^]� ���������̋A�������������U��j0�u�=  ��]���������������U��j0�u���  ��P�z=  ��]������U����E�j0�u�uP���  ��P�P=  ����M��@Q�@�Ѓ���]���������U����E�j0�u�u�uP��  ��P�=  ����M��@Q�@�Ѓ���]������U��j$�u��<  3Ƀ�������]�����U��j$�u�#�  ��P�<  3Ƀ�������]������������U����E�Sj$�u�uP��  ��P�<  ���3ۋI���I�E�P���у���[��]������������U����E�Sj$�u�u�uP�%�  ��P�,<  ���3ۋI���I�E�P���у���[��]���������U�졠��u�@�u���   j �Ѓ�]�U���u����u�@�u���   j �Ѓ�]��������������U�졠��@���  ]��������������U�졠��@0���   ]��������������U�졠����@0V���   W�u�M��uQ�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]��������������U���4���S�@V�u�@WV�С���M�@�����   3�SS�ЋM�E����S�@j���   �Ћ����M  3ɉM�d$ ��~k����M�@Q�@�С��j �@j��@�M�h��Q�С�����@�΋@<�Ћȡ��j��@j��@L�U�RQ���С���M�@Q�@�Ѓ����W�@0�u����   �M�Q�Ћ�����M܋@Q�@�С���M܋@Q�@W�С���M̋@Q�@�С�����@�΋@<�Ћȡ��j��@j��@L�U�RQ���С���M܋@Q�@�С���M�@�����   ��
j �MQ�MC�ЋM�E����A�Pj ���   Q�M�ҋ��������_��^[��]����U�졠��@0���   ]��������������U�졠��@0���   ]��������������U�졠��@0���   ]�������������̋�W��JR��A(�P$j j h����=  �������������̸�������������U���(V��W��M�Q���P(�V����t&���j �A0j ���   j j j j Wj jR�Ѓ�(����M�@Q�@�С���M�@Q�@�ЋN����t&���j �@0j ���   j �U�Rj jj?j Q�Ѓ�$����M�@Q�@�С���M�@Q�@�ЋN����u3��:����U�Rj j j h  
 j�U�R�E�    �@0h�  ���   jQ�Ћ}���(����M�@Q�@�Ѓ���u_3�^��]á���M�@Q�@�ЋN����t&���j �@0j ���   j �U�Rj j j8j Q�Ѓ�$����M�@Q�@�ЋN����t���j�@0Q�@P�Ѓ�����M�@Q�@�Ѓ��M��e���Ph   h  K j;�E�Ph	��h�  �����������M�@Q�@�Ѓ��M�臧���N��t���Q�@0�@X�Ѓ��N��t���Q�@0�@X�Ѓ��N��t&���j �@0j ���   j j j jj j jQ�Ѓ�(j�v$��5  ���   _^��]���U���V��Wj�N�\�  �F4    �F8    �F<    W��F(���h�   �@0�v�@�С���M�@Q�@�С��j �@j��@�M�h��Q�Ѓ��E�j j P�E�P���E��  �E�    �[�������M�@Q�@�Ѓ��Nj j��  _^��]������U���\���V�@W�@���M�Q�С��j �@j��@�M�h��Q���G(�Y������E��  �I�,��E�    �RP�E�P���   �Ћ�����I�E؋IP�ы���A�M؋@QV�С���M��@Q�@�С���M�@Q�@�С���M�@Q�@�M�Q�С����<�@�M�@<�Ћ��j��Qj��M�QP�BL�M���j j �E�P�E�P���&�������M�@Q�@�С���M؋@Q�@�С���Mȋ@Q�@�Ѓ��M�htats�ä�����j�@j�@0�M��С���G(�@���@,�$j�M��ЍE�P�E�P�E�P���E��  �E�    �_�������M����   Q� �Ѓ��4 tq����O0�@P�@h�ЋG4��t�w8�Ѓ��G<�G8    �G4    �/hh�hP	  hx�h  @�P  ���=�� t
�=�� t̡���O0�@P�@l�ЍM�����_^��]� ��U�졠���@�@V�@ W�}�����=MicMtc=ckhctG=fnic��   j�M�董���MP�أ���M����������M�@j�@4j��_�   ^��]� ����P���_��^��]� ���j �@hIicM���   ����=���uhtats�M��������j �@j�@0�M��ЍE�P�E�P�E�P���E��  �E�    �ط������M苀�   Q� �Ѓ��M��
����N�F   ��t���Q�@0�@�Ѓ��u��W�����_^��]� ��������U��mV��t3�^]� j�N��  j�L1  �N���F    ��t���Q�@0�@�Ѓ��   ^]� j�����  j�1  ��3�����������U���E�A(]� ��������������̍A�������������U��VW��~4 tU�I hh�h	  hx�h  @�GN  ���=�� t
�=�� t�j
�j=  ����v �@P�@�Ѓ���u_9F4u�����N0�@P�@h�Ѓ~4 tLhh�h5	  hx�h  @��M  ���=�� t
�=�� t̡���N0�@P�@l���K���_3�^]� �E�F8�E�F4���S�@P�N0�@l�Ѓ~4 t#j
��<  ����v �@P�@�Ѓ���u99F4uݡ���N0�@P�@h�Ћ~<�F<    ����N0�RP�Rl��[��_^]� [_3�^]� ���������U����M�V�q����M�����t �@4Q�@�Ѓ���t$��M�Q�u���R(�1�@0�u�@�Ћȃ���u�M�3�臠����^��]Ë�U�R�u�P �𡠴�M�@�@ �Ѓ��t����H0�E�IxP�u�у��M��>�����^��]��������U�졠�V�@j �u���   ��M�Ћ���u�    �F^]� ��u9Ft�   ^]� ���������U��V�uW��;uuz����M�@j ���   htsem�Ѕ�u\����M�@j ���   hrdem�Ѕ�u>�E�E�H��t1���j �@0�U�@,RVQ�Ѓ���t�u���r  _�   ^]� _3�^]� ���������������U�졠���@�@V�@W���M�Q�С���MЋ@Q�@�С�����@�MЋ��   Q�u�M�Q�M�Ћ�����I�E��IP�ы���A�M��@QV�С���M��@Q�@�С���M��@Q�@�M�Q�С���M��@Q�@�С���MЋ@Q�@�С�����@��@V�С���M��@V�@Q�Ѓ����  ����M��@Q�@�Ѓ�_^��]� ���������U���SV�u��;u��   ����M�@j ���   htsem�Ѕ���   ����M�@j ���   hrdem�Ѕ���   ����M�@Q�@�ЋM���E�P�E�P�u��E�    �X�����u3��4������@��@V�С���M�@V�@Q�Ѓ����  �   ����E�IP�I�у���^[��]� ^3�[��]� ���U������V�@�����   W��$�u��M���]�����u�E��    �F^��]� ��u�Ff.E����D{�   ^��]� ����U���SV�u��;u��   ����M�@j ���   htsem�Ѕ�um����M�@j ���   hrdem�Ѕ�uO�EW��H�E���t=���j �@0�U��@0RVQ�Ѓ���t!�E������$�|  ^�   [��]� ^3�[��]� �����U���0���V��W��M�Q�u�E��E��E��@�MЋ��   Q�M���~�~P�~H����uf�^f�V�    f�N^��]� ��u3�Ff.ß��Dz�Ff.��Dz�Ff.����D{�   ^��]� ��������U���4�ES�]V�uW�}�M�;�t;�t;���   ����M�@j ���   htsem�Ѕ���   ����M�@j ���   hrdem�Ѕ�ux�M�E��E��E�E�P�E�P�E�PW��E�P�E��E��E܉u�}�]��̺����t8�~E̋M�����f� �~E�f�@�~E�f�@�  �   _^[��]� _^3�[��]� �����U���0���V��W��E�����M�Q�u�E��@�MЋ��   Q�M���~ �~H�f�E�f�M���uf�F�    f�N^��]� ��u�E�P�FP��   ����t�   ^��]� ��������������U���SV�u��;u��   ����M�@j ���   htsem�Ѕ�u|����M�@j ���   hrdem�Ѕ�u^�M�E��E�P�uW��E�����E�P�E��u�������t,�~E���ċ�f� �~E�f�@�-  �   ^[��]� ^3�[��]� ������U���V�uW�}�f.���Dz�Ff.G���D{Y�G�Y����E��E��$�X> �F�]��Y�E��E��$�<> �E��]���f.E����D{_�   ^��]�_3�^��]����U��V��N�����t���Q�@0�@�Ѓ��E�F    t	V�)p������^]� ���������������U��V��~ �l�u����v�@4� �Ѓ��E�F    �F    t	V��o������^]� ��������U�����u�E�    �A]� ��u�A;Et�   ]� U�����u�E�    �A]� ��u�Af.E���D{�   ]� ����U�����u(�~Ef�A�~Ef�A�~E�    f�A]� ��u6�Af.E���Dz �Af.E���Dz�Af.E���D{�   ]� U��V�����u�~Ef�F�~E�    f�F^]� ��u�EP�FP��������t�   ^]� �U��V�����u �    ����P�FP�EP�B�Ѓ��"��u����M�@Q�@x�N�Ѕ�t�   ����M�@Q�@�Ѓ�^]� �������̡��Q�@L���   �Ѓ�������������U�졠��u�@L�u���   Q�Ѓ�]� ���������������U�졠�V�@L�񋀠   V�Ћȡ������u�@LQ�u���   V�Ѓ�^]� ���   �@P�Ћ��P���   �M�BH��^]� �������������̡��Q�@L��(  �Ѓ�������������U�졠��u�@L�u��,  Q�Ѓ�]� ��������������̡���@L� ������U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡���@L���   ��U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U�졠����@L�u�@Q�M�Q�ЋM��P�y����M�葔���E��]� ��������U�졠��u�@L�u�@Q�Ѓ�]� ��U�졠��u�@LQ���   �Ѓ�]� �̡��Q�@L�@�Ѓ���������������̡��Q�@L�@�Ѓ���������������̡��Q�@L�@�Ѓ����������������U���u����u�@L�u�@ Q�Ѓ�]� ���������������U�졠��u�@LQ��4  �Ѓ�]� ��U���u����u�@L�u�@$Q�Ѓ�]� ���������������U���u����u�@L�u�@(�uQ�Ѓ�]� �����������̡��Q�@L�@,�Ѓ���������������̡��Q�@L�@0�Ѓ���������������̡��Q�@L�@4�Ѓ���������������̡��j �@LQ�@8�Ѓ��������������U�졠��u�@L�u��  Q�Ѓ�]� ���������������U�졠��@L���   ]��������������U�졠��@L���   ]��������������U�졠��@L��l  ]��������������U�졠��@L���   ]��������������U�졠��@L���   ]��������������U�졠��@L���   ]��������������U�졠��@L���   ]��������������U�졠��@L���   ]��������������U�졠��@L���   ]��������������U�졠��u�@LQ�@<�Ѓ�]� �����U�졠��@L���   ]�������������̡��Q�@L�@��Y�U�졠��u�@L�u�@@Q�Ѓ�]� ��U�졠�j �@L�u�@DQ�Ѓ�]� ���U�졠�j�@L�u�@DQ�Ѓ�]� ���U�졠�j �@L�u�@HQ�Ѓ�]� ���U�졠�j�@L�u�@HQ�Ѓ�]� ��̡��Q�@L���   �Ѓ�������������U�졠����@L�u��  Q�M�Q�ЋM��P�����M������E��]� �����U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    觎  j �E�P�E�P���?  ���M�����  ��t3������M܋��   Q�@8�Ѓ�������E܋��   P�	�у���^[��]����������U���$V�E��P�M��E�   �E�   �E��  �E�    �E�    ��  j�E�P�E�P���?  �M���  ����M܋��   Q� �Ѓ�^��]�����U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    藍  j �E�P�E�P���v>  ���M����	�  ��t
�M�Mh��� ����M܋��   Q�@L�ЋM��P��h������E܋��   P�	�ыE��^[��]� ���������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    ��  j �E�P�E�P����=  ���M����Y�  ��t
�M�g��� ����M܋��   Q�@L�ЋM��P�+h������E܋��   P�	�ыE��^[��]� ���������U���$���V�u�E�    �E�    ���   ��@(�M�Q�Ѓ��E�P�M��E��  �E�    �E�    ��  j�E�P�E�P���=  �M�蕍  ����M܋��   Q� �Ѓ�^��]� ��������U���$���V�u�E�    �E�    ���   ��@(�M�Q�Ѓ��E�P�M��E��  �E�    �E�    莋  j�E�P�E�P���<  �M���  ����M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    ��  j �E�P�E�P����;  ���M���艌  ^��[tW��E��E������M܋��   Q�@<�Ѓ�����]��M܋��   Q� ���E�����]����������������U����EV�E��P�M�E�   �E��E��  �E�    �E�    �e�  j�E�P�EP���d;  �M�܋  ����M䋀�   Q� �Ѓ�^��]� ���������������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    ��  j �E�P�E�P����:  ���M����Y�  ��t3������M܋��   Q�@8�Ѓ�������E܋��   P�	�у���^[��]����������U���$�EV�E�E��P�M��E�   �E��  �E�    �E�    �I�  j�E�P�E�P���H:  �M����  ����M܋��   Q� �Ѓ�^��]� ���U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �׈  j �E�P�E�P���9  ���M����I�  ��t8����u���   W��	�����E�P�F�у���^[��]� ����M܋��   Q�@P���~ �u���f��~@���   �E܋	Pf�F�у���^[��]� ���U���$���V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    �އ  j�E�P�E�P����8  �M��U�  ����M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �g�  j �E�P�E�P���F8  ���M����و  ��t8����u���   W��	�����E�P�F�у���^[��]� ����M܋��   Q�@P���~ �u���f��~@���   �E܋	Pf�F�у���^[��]� ���U���$���V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    �n�  j�E�P�E�P���m7  �M���  ����M܋��   Q� �Ѓ�^��]� ��������U�졠����@Lj�u���   Q�M�Q�ЋM�~ f��~@��f�A����]� U�졠����@Lj �u���   Q�M�Q�ЋM�~ f��~@��f�A����]� U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �w�  j �E�P�E�P���V6  ���M�����  ��t8����u���   W��	�����E�P�F�у���^[��]� ����M܋��   Q�@P���~ �u���f��~@���   �E܋	Pf�F�у���^[��]� ���U���$���V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    �~�  j�E�P�E�P���}5  �M����  ����M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    ��  j �E�P�E�P����4  ���M����y�  ��t8����u���   W��	�����E�P�F�у���^[��]� ����M܋��   Q�@P���~ �u���f��~@���   �E܋	Pf�F�у���^[��]� ���U���$���V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    ��  j�E�P�E�P���4  �M�腄  ����M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    藂  j �E�P�E�P���v3  ���M����	�  ��t3������M܋��   Q�@8�Ѓ�������E܋��   P�	�у���^[��]����������U���$�EV�E�E��P�M��E�   �E��  �E�    �E�    ���  j�E�P�E�P����2  �M��p�  ����M܋��   Q� �Ѓ�^��]� ���U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    臁  j �E�P�E�P���f2  ���M������  ��t8����u���   W��	�����E�P�F�у���^[��]� ����M܋��   Q�@P���~ �u���f��~@���   �E܋	Pf�F�у���^[��]� ���U���$���V�u�E�    �E�    ���   ��@,�M�Q�Ѓ��E�P�M��E��  �E�    �E�    莀  j�E�P�E�P���1  �M���  ����M܋��   Q� �Ѓ�^��]� ��������U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    ��  j �E�P�E�P����0  ���M���艁  ��t3������M܋��   Q�@8�Ѓ�������E܋��   P�	�у���^[��]����������U���$�EV�E�E��P�M��E�   �E��  �E�    �E�    �y  j�E�P�E�P���x0  �M����  ����M܋��   Q� �Ѓ�^��]� ���U���$SV�E��P�M��E�    �E�    �E��  �E�    �E�    �  j �E�P�E�P����/  ���M����y�  ��t3������M܋��   Q�@8�Ѓ�������E܋��   P�	�у���^[��]����������U���$�EV�E�E��P�M��E�   �E��  �E�    �E�    �i~  h�   �E�P�E�P���e/  �M���  ����M܋��   Q� �Ѓ�^��]� �������t��t��t3�ø   ���̡��Q�@L�@L�Ѓ���������������̡��Q�@L�@P�Ѓ����������������U���u����u�@L�u���  Q�Ѓ�]� ������������U�졠��u�@LQ��  �Ѓ�]� ��U�졠��u�@LQ���   �Ѓ�]� �̡��Q�@L�@X�Ѓ����������������U���u����u�@L�u�@\Q�Ѓ�]� ���������������U�졠���0�@LS�@V���Ћ؅�u^[��]� W�M��}���u�E�Eء���E�    �E�    �E�    �E�    �E�    �]Ћ@h]  �@0�M��С��j ���   j �@S���Ѕ���   ���S�@L�@�Ћ�������   �d$ ������   �΋R(�ҋ��E�Ph�   �u���  ����tq�M��tj���j ���   ���   �ЋЅ�tO���V���   �ʋ@<�С���M苀�   Q���   �Ѓ���t���V�@@�@�Ѓ������d����*���S�@@�@�С���M苀�   Q���   �Ѓ�3ۍM��0  �M��|��_^��[��]� ������������̡��Q�@L�@`�Ѓ���������������̡��Q�@L�@d�Ѓ����������������U�졠��u�@LQ�@h�Ѓ�]� ����̡��Q�@L��D  �Ѓ������������̡��Q�@L�@l�Ѓ����������������U�졠��u�@LQ���   �Ѓ�]� �̡���@L�@�����U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��Q�@L���   ��Y�������������̡��Q�@L���   �Ѓ�������������U���u����u�@L�u���   �u�uQ�Ѓ�]� ������U���u����u�@L�u���   Q�Ѓ�]� ������������U���u����u�@L�u��   �uQ�Ѓ�]� ���������U���u����u�@L�u��   Q�Ѓ�]� ������������U�졠��@L��H  ]�������������̡���@L��L  ��U�졠��@L��P  ]��������������U�졠��@L��T  ]��������������U�졠��@L��p  ]��������������U�졠��@L��t  ]��������������U�졠��@L���  ]��������������U�졠��@L���  ]��������������U�졠��@L���  ]�������������̡���@L���  �ࡠ��@L���  ��U��U$V�u�Eh�h�h�h�R�u �q�u�Q�u������@L�$�u���   VQ�Ѓ�4^]�  �������̡���@���   �ࡠ��@���   ��U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠�V�@�u���   �6�Ѓ��    ^]������������U�졠�V�@L�@�Ћ���u^]��u���j �u�@�u���  �uV�Ѓ���u���V�@@�@�Ѓ�3���^]���������U���u���j �H�u�E�� P�u���  �u�Ѓ�]����U�졠��@���   ]��������������U�졠��@L���   ]��������������U���u(����u �@�u���  �u�u�u�u�u$�u�Ѓ�$]��������������U�졠�V�u0�p�u,�E����P�Q���u���  �u�Ѓ�,�M���Q����^]�U�졠��@���  ]��������������U��� ����E�    �E�    �E�    �E�    �E�    �E�    �E�    ���   V���   �Ћu�E���t8��t4���j�QLP���   ���ЋE��E�E�Ph=���u���
  ������   ����M����   Q���   �Ѓ��M��E�    �  ��^��]���������������U��� ����E�    �E�    �E�    �E�    �E�    �E�    �E�    ���   V���   �Ћu�E���t8��t4���j�QLP���   ���ЋE��E�E�Ph<���u��*
  ������   ����M����   Q���   �Ѓ��M��E�    ��   ��^��]���������������U�졠��@L���   ]��������������U�졠��@L���   ]�������������̡���@L��  �ࡠ��@L��@  ��U��M�]� �����U��M�u��P]�U��M�u��u�P]��������������U���u�M�u��u�u�P]�������̡�����   �AP���   ��Y��������U�졠��u�@8Q�@D�Ѓ�]� ����̡���@8�@<�����U�졠�V�@8�u�@@�6�Ѓ��    ^]���������������U���u����u�@8�u�@�u�u�uQ�Ѓ�]� ������U���u����u�@8�u�@�u�uQ�Ѓ�]� ��������̡���@8� ������U�졠�V�@8�u�@�6�Ѓ��    ^]���������������U���u����u�@8�u�@Q�Ѓ�]� ���������������U�졠��u�@8�u�@Q�Ѓ�]� �̡��Q�@8�@�Ѓ����������������U�졠��u�@8Q�@ �Ѓ�]� �����U���u����u�@8�u�@$�u�uQ�Ѓ�]� ���������U�졠��u�@8�u�@(Q�Ѓ�]� ��U���u����u�@8�u�@,Q�Ѓ�]� ���������������U���u����u�@8�u�@Q�Ѓ�]� ���������������U�졠��u�@8�u�@0Q�Ѓ�]� ��U���u����u�@8�u�@4Q�Ѓ�]� ���������������U�졠��u�@8Q�@8�Ѓ�]� �����U��M����P�APP�A@P�A0P�A P�AP���   Q�u�Ѓ�]�������������̡���@���   �ࡠ��@���  ��U�졠��@�@,]�����������������U�졠��@���  ]��������������U�졠�V�H�u�IV�ы��V�I�I8�у���^]����̡���@�@<�����U�졠��@���  ]��������������U�졠��@�@@]����������������̡���@�@D����̡���@�@H�����U�졠��@�@L]�����������������U�졠��@�@P]�����������������U�졠��@��<  ]��������������U�졠��@��,  ]��������������U���u����u�@�u���   �u�uh�:  �Ѓ�]�����U�졠��@�@]�����������������U�졠��� �@�M��@Q�С��j �@j��@�M�hT�Q�С���M��@Q�@�С���M��@Q�@�M�Q�С���� �@�M��@<�Ћ��j��Qj��u�M�P�BL�С���M��@Q�@�С���M��@Q�@�С���M��@Q�@�Ѓ���]����U�졠��@���  ]��������������U�졠��@��8  ]��������������U�졠����@V��  �M�WQ�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]����U�졠����@V��  �M�WQ�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]����U�졠��@��x  ]��������������U�졠��@��|  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@�@T]�����������������U�졠��@�@X]�����������������U�졠��@�@\]����������������̡���@�@`�����U�졠��@���  ]�������������̡���@�@d����̡���@�@h�����U�졠��@�@l]�����������������U�졠��@�@p]����������������̡���@���  ��U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@�@t]�����������������U�졠��@��D  ]��������������U�졠��@��  ]��������������U�졠��@�@x]�����������������U�졠��@��@  ]��������������U��V�u����D�����V�I�u�I|�у���^]���������U�졠��@���   ]��������������U�졠��@���  ]��������������U�졠��@��h  ]��������������U�졠��@���  ]�������������̡���@���   ��U��V�u���"j�����V�I���   �у���^]��������̡���@��`  �ࡠ��@���  ��U�졠��@��  ]��������������U�졠����@�u���   �M�Q�ЋM�~ f��~@f�A�~@��f�A����]������������U�졠��@���  ]��������������U���u�E������@�D$�E���   �$�u�Ѓ�]�����������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@��   ]��������������U�졠��@��  ]��������������U�졠��@��l  ]�������������̡���@���  ��U�졠��@���  ]��������������U�졠����@�u���  �u�M�Q�ЋM��P�B���M���B���E��]������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠����@V���  W�u�M�Q�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]�U�졠����@V���  W�u�M�Q�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]�U�졠��@���  ]��������������U�졠��@���  ]��������������U�������U��@R���   �U�R�U�RQ�Ѓ����#E���]����������������U�������U��@R���   �U�R�U�RQ�Ѓ����#E���]����������������U�������U��@R���   �U�R�U�RQ�Ѓ����#E���]����������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@���   ]��������������U�졠��@��  ]��������������U�졠��@��\  ]��������������U�졠����H�u��t  �u�E�P�у�����?���M��N?���E��]��������U�졠��@��H  ]��������������U�졠��@��T  ]�������������̡���@��p  ��U�졠��@��8  ]��������������U���  �H�3ŉE��EP�u������h   P�
 ����x	=�  |5�/h�hR  hx�h  @�  ���=�� t
�=�� t��E� ����������@Q��4  hX��ЋM�3̓��f�  ��]����������������������U���u(�E�u$�P�u ����u�@0�u���   �u�u�uRQ�Ѓ�(]�$ ������U���u(�E�u$�P�u ����u�@0�u���   �u�u�uRQ�Ѓ�(]�$ ������U���u(����u$�@0�u ���   �u�u�u�u�u�uQ�Ѓ�(]�$ ���������̡��Q�@0���   �Ѓ�������������U�졠��u�@0�u���   Q�Ѓ�]� ���������������U���u����u�@0�u���   �uQ�Ѓ�]� ��������̡��Q�@0���   �Ѓ�������������U���u����u�@0�u���   �uQ�Ѓ�]� ��������̡���@0���   ��U�졠�V�@0�u���   �6�Ѓ��    ^]������������U�졠����@V�u��X  �u�M��uQ�Ћuj �    �F    ���P���   V�I�ы���E����   P�	�у� ��^��]����������U�졠����@V���  W�u�M�Q�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]�U���4VhLGOg�M��`�����j �IP�E�hicMCP��X  �Ћ�����E�    �E�    ���   j �@R�M�Q�С���M����   Q� �Ѓ� �M��i`������M����   Q�@T�Ѓ���u
�M��_��� ����M����   Q�@T�ЋM��P�`������E����   P�	�ыE��^��]������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠����@V��t  Wj �u�M��u�u�uQ�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у�(��_^��]������U�졠����@V�u���  �u�M��u�uQ�Ћuj �    �F    ���P���   V�I�ы���E����   P�	�у�$��^��]�������U�졠���4�@��p  �Ѕ���   h���M��U^������u�@h���@4�M��С���u�@h���@4�M��С��j �@�M̋�X  Q�M�hicMCQ�Ћ�����E�    �E�    ���   j �@R�M�Q�С���M����   Q� �С���M����   Q� �Ѓ�$�M���]����]����������U�졠���4�@V��p  �Ѕ�u����u�HV�I�у���^��]�Wh!���M��\]������u�@h!���@4�M��С��j �@�M̋�X  Q�M�hicMCQ�Ћ�����E�    �E�    ���   j �@R�M�Q�С���M����   Q� �С���M����   Q�@H�Ћ���}�IW�I���ы��W�AV�@�Ћ���E����   P�	�у�4�M���\����_^��]������������U�졠���4�@V��p  �Ѕ�u����u�HV�I�у���^��]�Wh����M��<\������u�@h����@4�M��С��j �@�M̋�X  Q�M�hicMCQ�Ћ�����E�    �E�    ���   j �@R�M�Q�С���M����   Q� �С���M����   Q�@H�Ћ���}�IW�I���ы��W�AV�@�Ћ���E����   P�	�у�4�M��[����_^��]������������U�졠���4�@��p  �Ѕ�u��]�Vh#���M��4[������u�@h#���@4�M��С��j �@�M̋�X  Q�M�hicMCQ�Ћ�����E�    �E�    ���   j �@R�M�Q�С���M����   Q� �С���M����   Q�@8�Ћ�������   �E��	P�у�(�M���Z����^��]�������U�졠���4�@��p  �Ѕ�u��]�Vhs���M��TZ������u�@hs���@4�M��С��j �@�M̋�X  Q�M�hicMCQ�Ћ�����E�    �E�    ���   j �@R�M�Q�С���M����   Q� �С���M����   Q�@8�Ћ�������   �E��	P�у�(�M���Y����^��]������̡���@��d  ��U�졠��@��h  ]��������������U�졠��@��l  ]��������������U�졠��@���  ]�������������̡���@���  ��U�졠��@���  ]��������������U�졠��@��   ]�������������̡���@��P  �ࡠ��@���  ��U�졠����@�u���  �M�Q�ЋM��P�X���M���X���E��]���������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@��l  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@��$  ]��������������U�졠��@��(  ]��������������U�졠��@��,  ]�������������̡���@��0  �ࡠ��@��<  ��U�졠��@��  ]��������������U�졠��@��`  ]��������������U�졠��@��\  ]��������������U��� V����u3�^��]�W�v�v�v�v�}  ����u_^��]������E�Pjd�E�P�E�   �E�觀  Pjd���m�  ����M����   Q� �С���M����   Q� �Ѓ���_^��]�������������U���V��> u3�^��]�SW��   �΋��{  ��褀  �E�����   j jSW���l}  ����   ��<  ��t�M�j j��~  �N�V�C�P�G�P�Fj Hj �P�FH�PQ�R�u���}  ����M��E�Pjd�E�   �E��~  ����M싀�   Q� �ЋE���_[^��]ÍE�P��  ��3�_[^��]����������U���(V����u�F^��]�����E�Pjd�E�P�E�   �E��6  ���P���   �@<���]�����M؋��   Q� �С���M苀�   Q� ���M��N��f. ����D{fn�����^��,ȋ�^��]������������U���(V����u�F^��]�����E�Pjd�E�P�E�   �E��~  ���P���   �@<���]�����M؋��   Q� �С���M苀�   Q� ���M��N��f. ����D{fn�����^��,ȋ�^��]������������U��E���� ]��U����S�]#ètc��th���
��th��hX��^������uhX��N�������   @t�u�u�(  ����    uh��hX�������[]���������U���  �H�3ŉE�����M�    �   E�S�]���#è��   �EPQ������h�  P��  ����th���
��th��hX�������������PhX���������   @t�u�u�b   ����    uh��hX��X������M�3�[�G�  ��]������������������U��]���  �������U��]��  �������U���L  �H�3ŉE�V�u������P�^�  ������P��  Ph���E�j?P��  �u�E�VPh��������h�  P�2   ������PhX������M���83�^��  ��]����������������U��V�u��3�^]�W�}�EP�uVW�/�  ����x;�|l�D7� _�F�^]����t<h��hX��/���hx�hX�� ���h��j+����h��hX������� �=�� t
�=�� t��D7� �F�_^]�����A    �    �A    �A   �����U���u����u�@@�u�@Q�Ѓ�]� ���������������U�졠��u�@@Q�@�Ѓ�]� �����U�졠��u�@@�u�@Q�Ѓ�]� ��U�졠��u�@@Q�@ �Ѓ�]� �����U�졠����   �@]��������������U�졠����   �@]��������������U�졠����   �@ ]�������������̡�����   �@$��U�졠����   ���   ]�����������U�졠����   ��D  ]�����������U�졠��u�@@Q�@L�Ѓ�]� ����̡��Q�@@�@H�Ѓ����������������U�졠����   ���   ]�����������U�졠����   ���   ]����������̡��Q�@H���   �Ѓ�������������U��V��M��t2�U������   ��t�@@R��^]� �U�@D��tR��^]� V��^]� �����������̡���@@�@0�����U��V�u���t���Q�@@�@�Ѓ��    ^]����������U�졠�V�@@��@V�ЋЋE����t��#��С��R�@@V�@�Ѓ�^]� �U���u �E��������   �$�u���   �u�u�u��]� ����������U�졠����   ���   ]����������̡��Q�@H���   �Ѓ�������������U�졠��u�@HQ��d  �Ѓ�]� �̡���@@�@T�����U�졠��@@�@X]�����������������U�졠��@@�@\]����������������̡���@@�@`�����U�졠��@@�@d]�����������������U�졠��@@�@h]�����������������U�졠��@@�@l]�����������������U�졠��@@���   ]�������������̡���@@�@t����̡���@@�@x�����U�졠��@@�@|]����������������̡���@@���   ��U�졠��@@���   ]�������������̡���@@���   �ࡠ����   �@t��U�졠��@@���   ]��������������U�졠��@@���   ]��������������U�졠��@@���   ]��������������U�졠��@@���   ]��������������U�졠��@@���   ]��������������U�졠��@@���   ]��������������U�졠��@@���   ]��������������U��V�u���t���Q�@@�@�Ѓ��    ^]���������̡���@@�@0�����U�졠�j�@@�M�@4Qj �Ѓ�]����U�졠�j�@@�M�@4Qh   @�Ѓ�]�U�졠��u�@@�u�@4j �Ѓ�]���̡���@|� ������U��V�u���t���Q�@|�@�Ѓ��    ^]���������̡���@|�@ �����U��V�u���t���Q�@|�@(�Ѓ��    ^]����������U�졠��@ �@H]�����������������U��}qF uGW�}��t>����u���   �ϋ@D�С���u�@@�@,�Ћ�����ЋAW�u�@p����_]������������U�졠��@��T  ]��������������U�졠�S�@@V�@,W�u�Ћ���u�I@�؋I,�ы�����yh��hE  �ˋ��8J��Ph��hE  ���&J��P��T  �Ѓ�_^[]������U��E�+u&�Q+Pu�Q+Pu�Q+Pu�Q+Pu�Q+P3�����]� ���U��E�+u&�Q+Pu�Q+Pu�Q+Pu�Q+Pu�Q+P3�����]� ���U��E�+u&�Q+Pu�Q+Pu�Q+Pu�Q+Pu�Q+P3�����]� ���U��E�+u&�Q+Pu�Q+Pu�Q+Pu�Q+Pu�Q+P3�����]� ���U��E�+u&�Q+Pu�Q+Pu�Q+Pu�Q+Pu�Q+P3�����]� ���U��E�+u&�Q+Pu�Q+Pu�Q+Pu�Q+Pu�Q+P3�����]� ���U��E�M�+t��]ËP+Qu�P+Qu�P+Qu�P+Qu܋@+A]������U���Vh��h�   h�f ����  ����t:���   ��t0�M�Q���ЋM�~ f��~@f�A�~@f�A��^��]� �E^� �  �@   �@   �@    �@    �@    ��]� ���������������U��Vh��h�   h�f ���v�  ����t���   ��t�u���u�u��^]� ���h��h�   h�f �<�  ����t���   ��t��3��������U��h��h�   h�f �	�  ����t���   ��t]��]����U���Vh��h�   h�f ���ӏ  ����t:���   ��t0�M�Q���ЋM�~ f��~@f�A�~@f�A��^��]� �E^� �  �@   �@   �@    �@    �@    ��]� ���������������U��Vh��h�   h�f ���6�  ����t���   ��t�u���u�u��^]� ���U��Qh��h�   h�f ���  ����t���   �E���t�u�U�����]������]��������������U���h��h�   h�f 覎  ����tE���   ��t;�E���M��$Q�ЋM�~ f��~@f�A�~@��f�A����]ËE� �  �@   �@   �@    �@    �@    ��]�����������U��h��h�   h�f �	�  ����t���   ��t]��]����U���h��h�   h�f �E��  �E�   �E�   �E�    �E�    �E�    謍  ����t���   ��t	�M�Q�Ѓ�h��h�   h�f �~�  ����t���   ��t�u�M�Q�Ѓ���]ËE�~E�f� �~E�f�@�~E�f�@��]����������U��h��h�   h�f ��  ����t���   ��t]���M�E�~f� �~Af�@�~Af�@3�]����������������U��h��h�   h�f 蹌  ����t���   ��t]���M�E�~f� �~Af�@�~Af�@3�]����������������U��h��h�   h�f �Y�  ����t���   ��t]��3�]��U���Vh��h�   h�f �%�  ����tX���   ��tNW�u�M��uQ�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]á���u�HV�I�у���^��]������������U��VWh��h�   h�f 臋  ������tI���    t@�u ����u�@�u�@����V�С���M�@V�@Q�Ћ��   ���Ѓ����3�����E�IP�I�у���_^]���������U��VWh��h�   h�f ���  ������tI���    t@�u ����u�@�u�@����V�С���M�@V�@Q�Ћ��   ���Ѓ����3�����E�IP�I�у���_^]���������U���Vh��h�   h�f �e�  ����tX���   ��tNW�u�M��uQ�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]á���u�HV�I�у���^��]������������U���Vh��h�   h�f �ŉ  ����tU���   ��tKW�u�M�Q�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]á���u�HV�I�у���^��]���������������U���Vh��h�   h�f �%�  ����tU���   ��tKW�u�M�Q�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]á���u�HV�I�у���^��]���������������U��h��h�   h�f 艈  ����t���   ��t]��]����U��h��h�   h�f �Y�  ����t���   ��t]��]����U��h���uh�f �+�  ��]�������U�졠��@ �@h]�����������������U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U�졠��u�@ Q�@�Ѓ�]� �����U�졠��u�@ Q�@�Ѓ�]� ����̡��Q�@ �@��Y�U��VW�}����?=�����W�J V�I�у���_^]� ����U�졠��u�@ Q�@ �Ѓ�]� ����̡��Q�@ �@,�Ѓ���������������̡��Q�@ �@0�Ѓ����������������U�졠��u�@ Q�@4�Ѓ�]� ����̡���@ � ������U��V�u���t���Q�@ �@�Ѓ��    ^]����������U�졠��u�@T�u�@Q�Ѓ�]� ��U�졠��u�@TQ�@�Ѓ�]� �����U�졠��u�@TQ�@�Ѓ�]� �����U�졠����@T�u�@<Q�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� �����������U�졠��@T� ]��U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��hG  �@T� �Ѓ�������������U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U�졠�Q�u�@H�u���  �u�Ѓ�]� ������������U�졠��E�@H���@�$Q�Ѓ�]� ����������̡��j �@HQ���   �Ѓ�����������U�졠��u�@Hj ���   Q�Ѓ�]� ���j�@HQ���   �Ѓ�����������U�졠��u�@Hj���   Q�Ѓ�]� ���j�@HQ���   �Ѓ����������U�졠��u�@Hj���   Q�Ѓ�]� ���Q�@H���  �Ѓ�������������U�졠��u�@HQ���  �Ѓ�]� ��U�졠��u�@HQ���  �Ѓ�]� ��U�졠��u�@HQ���  �Ѓ�]� ��U�졠��u�@H�u��  Q�Ѓ�]� ���������������U�졠��u�@H�u��  Q�Ѓ�]� ��������������̡��Q�@H���   �Ѓ�������������U��VW�u���!.  ������t����u�AHV���   W�Ѓ���_^]� �������U��VW�u���u�.  ������t����u�AHV���   W�Ѓ���_^]� ����U�졠��u�@H�u���   Q�Ѓ�]� ���������������U�졠��u�@H�u���   Q�Ѓ�]� ���������������U�졠��u�@HQ���   �Ѓ�]� �̡��Q�@H���  �Ѓ�������������U���u����u�@H�u���  �u�uQ�Ѓ�]� ������U�졠����@HS���   Vj ��h�  V�   �Ћȃ���t8���Q�@@�@,�Ћȃ���u^[��]� ���j�@h�  ���   �Ћ؋��j �IHh�  ���   V�у��} u^�   [��]� Wh�  �>,  ��������   ���j �IHW���   V�у��M���6������u�@h�  �@0�M��С���E�@���@,�$h�  �M��С��S�@h�  �@0�M��С��j�@@�M�@(QW�Ѓ��M���6��_^�   [��]� _^3�[��]� ��������̡��Q�@H���   ��Y��������������U�졠��u�@HQ���  �Ѓ�]� ��U�졠��u�@HQ���  �Ѓ�]� �̡��Q�@H��4  �Ѓ�������������U�졠��@H� ]��U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U��S�]V�uW�> ��u3���S�@HW���   �Ѓ���u���j�@HW���   �Ѓ���t�   ��u����   ���W�@H���   �Ѓ��} u!�u����u�@H�u���  VSW�Ѓ��I�ΉM��t@�u��u���V�u�@HQ���  SW�С���M���   ���@(�ЋȉE��uǋu�E�8 u���W�@H���   �Ѓ���t3���   �EW�����@H��u$���   �С��S�@HW���   �Ѓ�_^[]� ���   �С�����} �@Hu�u���  j �uVSW�Ѓ�_^[]� � h  �Ѓ��E��u_^[]� ����΋��   �@x�Ћ��P���   �M�B|�Ѕ�tP�u���j �u�@HV���  SW�Ћȃ���t����u���   �@H�С���΋��   �@(�Ћ���u��E_^[]� U���u����u�@H�u���  �u�uQ�Ѓ�]� �����̡��Q�@H���   ��Y�������������̡��Q�@H���   �Ѓ�������������U�졠��u�@H�u���   Q�Ѓ�]� ��������������̡��Q�@H���   ��Y�������������̡��Q�@H��t  ��Y�������������̡��Q�@H��P  �Ѓ������������̡��Q�@H��T  �Ѓ������������̡��Q�@H��X  �Ѓ�������������U�졠����@HQ��\  �M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ����������̡��Q�@H��`  �Ѓ�������������U�졠��u�@HQ��d  �Ѓ�]� ��U�졠��E�@H����h  �$Q�Ѓ�]� ��������U�졠��E�@H����t  �$Q�Ѓ�]� ��������U�졠��E�@H����l  �$Q�Ѓ�]� ��������U�졠��u�@HQ��p  �Ѓ�]� ��U���u����u�@H�u���  �uQ�Ѓ�]� ���������U���u����u�@H�u���  �u�u�uQ�Ѓ�]� ��̡��h�  �@H� �Ѓ�������������U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��Q�@H���   �Ѓ������������̡��Q�@H���   �Ѓ�������������U�졠��u�@HQ���   �Ѓ�]� ��U�졠��u�@HQ���   �Ѓ�]� ��U�졠��u�@H�u���  Q�Ѓ�]� ���������������U�졠��u�@H�u��   Q�Ѓ�]� ���������������U���u����E�@H�����  �$Q�Ѓ�]� �����U�졠�V�@Hh  � �Ћ�������   �uh�  �%  �Ѓ���t^���j �AHR���   V���uh(  ��$  �Ѓ���t3���j �AHR���   V�С�������   j �@j���Ћ�^]á��V�@@�@�Ѓ�3�^]�����U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��Q�@H��  �Ѓ������������̡��Q�@H��  �Ѓ������������̡��Q�@H���  �Ѓ������������̡��Q�@H���  �Ѓ������������̡��Q�@H���  �Ѓ�������������U�졠��u�@H�u��  Q�Ѓ�]� ���������������U���u����u�@H�u��   Q�Ѓ�]� ������������U���u����u�@H�u��|  �uQ�Ѓ�]� ���������U��EV���u����@H���  �'��u����@H���  ���u(����@H���  V�Ѓ���tP�u���   ^]� 3�^]� ����������U���SW���!  �؅���   �} ��   ���V�AHj ��p  h�  W�Ћ�����IHh�  ���   W�u��������E����   �u3��Ή}���  ����   �E�P�E�P�u��W�  ��t\�u�;u�T������u�U����ɋD�;D�t-����Hl����P�E�p�A�ЋD������tP���  F;u�~��}��MG�}��`  �u;��v���^_��[��]� _3�[��]� U������V�@Hj ��p  ��h�  V�u��Ѓ��E���u^��]� �EW��u����@H���  �+��u����@H���  ����T  ����@H���  V�Ћ������6  S���/  ���h�  �@H3ۋ��   V�]��Ѓ�����   �E����s�E����M�@lS�q�@�Ћ؃�����   ����s�I\�u�I,�у���t�F�P���V  ����s�@\�u�@,�Ѓ���t�F�P���1  �M�;At"����s�@\�u�@,�Ѓ���tV���  ����s�@\�u�@,�Ѓ���t�FP����  ����]��@H�E���   h�  �u�C�]����Ѓ�;�����[_�   ^��]� _3�^��]� ������̡��Q�@H���  �Ѓ�������������U�졠��u�@H�u���  Q�Ѓ�]� ���������������U���u����u�@H�u���  Q�Ѓ�]� �����������̡��Q�@H���  �Ѓ������������̡��Q�@H���  �Ѓ�������������U�졠��u�@HQ��  �Ѓ�]� ��U�졠��u�@HQ��  �Ѓ�]� �̡��Q�@H��  �Ѓ�������������U�졠��u�@HQ��  �Ѓ�]� �̡��Q�@H��T  �Ѓ�������������U�졠��u�@H�u��  Q�Ѓ�]� ���������������U�졠��u�@HQ��8  �Ѓ�]� ��U�졠��u�@HQ��<  �Ѓ�]� ��U���u����u�@H�u��@  Q�Ѓ�]� ������������U�졠��u�@HQ���  �Ѓ�]� ��U�졠��u�@HQ��H  �Ѓ�]� �̡��Q�@H��L  ��Y��������������U�졠�V�@Hh�  � �Ћ�����u^]á���u�@H�u��  V�Ѓ���u���V�@@�@�Ѓ�3���^]����������U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U���u����u�@H�u��   Q�Ѓ�]� ������������U�졠��E�@H����$  �$Q�Ѓ�]� �������̡��Q�@H��(  �Ѓ�������������U�졠��u�@H�u��,  Q�Ѓ�]� ��������������̡���@H��  ��U�졠��@H��  ]�������������̡��V�@@��@,WV�Ћ�����ȋBj ���   h�  �Ћ��h�  �IHV���   ���у���
��t_3�^Ë�_^�̡��Q�@@�@,�Ћ�����ЋAj ���   h�  �������U�졠��E�@H����  �u�u���$Q�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ��������U�졠��E�@H����  �u�u���$Q�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� �������̡��Q�@H���  �Ѓ�������������U�졠��u�@H�u��8  Q�Ѓ�]� ���������������U���u����E�@H����0  �$�uQ�Ѓ�]� ��U�졠��@H�@]�����������������U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U���u �E�u������@H�$�u���   �u�u�Ѓ�]�������������U���u�E������@H�$�u���   �u�u�Ѓ�]�����������������    ���������̡��j�@H�1��|  �Ѓ����������U�졠�V�@H�u��x  ����3Ƀ������^��]� ���̡��j �@H�1��|  �Ѓ����������U��fnE�M����YE�X@��,�;�}��]�;EOE]����������������U���L���S�@HV�u���   Wh�  V�Ћ��3��IHW���   h�  V�E���3ۃ��E��}��}�]�9]���
  ����΋��   �@��=�  ����>  �@HS���   h:  V�Ћ��h�  �IHV���   �E��ы��S�IHh�  ���   V�E܉]��ы���u�IH����  �u��ы���u�IH�Eċ��  �у�(�E�9]�~y�^3��Eą�tSj�V���J�  ���tD�M��@�|� ���M�~�� ��%�������;�u+�Ȁ  �M�;�OȉM��M�腀  ���;Cu�����F��;u�|�3ۋu�����   j �u����  ����  ���  ��ty���v  �M�;�uk����ȋ�����������E��M��Uș;�u9U�uh��h�  Q��������3��E�����  �M��:  �M�I��QP�u��Ǧ  ���E왋ȋ�����������E��M��Uș;�u9U�uh��h�  Q�h������3��E���  �E�@��P�u��u��a�  �E�����~A����ȋ��������;�u;�uh��h�  Q�-������؉E��3ۉ]����  ����u�@Hj���  WV�Ѓ�����  �}���t jV���  ���{  ���T  ���E��3��}ࡠ�j �@Hh�  ���   V��3�3҃��E�U��M�9M��  �u���u���]�Eą��&  j�Q����  ����  �M��@�|� ���M�~�� ��%�������9E���  �9~  �E��E�3�3��E�    9p~h�I ��������ШtL�U�������������������L��B�D��A�D��B�D��A�D��B�D��A�D����E�G;x|����  �ƙ+�����~SPS�M��  �U��M�R3ۍ<��E�+��E��}ԋÐ;E��  �}� �E�����E��M�t:�I�M��~��M�f�9�}��~D��}�f�D9�M��~D��E��M�f�D8�I�M��~�f��~D�f�G�~D��M�f�G;�}w�}�����    9O�uc�����������w>�$��x�M�U�����-�M�U���T���M�U���T���M�U���T���U��M؃���;�|��}ԋE�B��@�U��}ԉE�;������;E��  �u��  �U��3�;F�Ã}� �]���   �R�ǋF��}��@�~�f��~D�f�A�~D�f�A�F��@�~�f�A�~D�f�A �~D�f�A(��ϋ}��@�~����Rf�D�0�~Af�D�8�~Af�D�@��t0�F�M��@�~����Rf�D�H�~Af�D�P�~Af�D�X�F��]�}�@�~ǍǍRf���~Af�D��~A��f�D��F��V��@B�~ǍǍRf���~Af�D��~A��f�D���V�B�@�~ǍǍRf���~Af�D��~A�ˋ]�f�D��B�U���t8�F�]�@�~ǍǍRf���~Af�D��~Af�D��VB�U����F��uȋU��M̋}�A���M̉u�;M�������E�E��E�P�����E��E��E�P�������c  �]�E�P�]������E��E��E�P�����E�E��E�P�s�����3�_^[��]Ë��   �΋@��=  �  ���j �@Hh(  ���   V�Ћ��h(  �IHV���   �E��ы؃�3��]ą���  ~"�U���    ��t�|� �<Ou���@;�|�E왋ȋ�����������E��M��U��;�u9U�uh��h~  Q�K��������3ɉM�M���tg�E�@��P�u�Q�E�  �Ù�ȋ����������;�u;�uh��h�  Q��������ȉE��3ɉM�M���u�E�E��E�P�4�����_^3�[��]Í�    P�u�Q�ן  ����]�IH�ǋ�   �+���PWS�E��у���u�E�P��  �E�P��  ��3�_^[��]Ë��ڬ���ˉE��  �M�3�3�3����}̉]��u�9U��-  �I ��    �E�����  3����|   �M��R�w���[�]�Ë]����    �~ f��~@f�A�~@f�A�~@f�A�~@ f�A �~@(f�A(��0�MȋM�F��G;4�Mȍ@|��]��u��M�|� ��    tj�M��}��@�~����RBf���~Af�D��~A�M�f�D��[�~����RBf���~Af�D��~A�M�f�D���    �]�F�u�;u�������}̋U�3���~!���$    �d$ �D�    ��   @;�|�E�P�M��@������E�E��E�P�.������   _^[��]ÍI �r�r�r�r������������U���u�E������@H�$�u���  �u�Ѓ�]���U�졠��@H���  ]��������������U�졠��@H���  ]��������������U���u0�E(������@H�$�u$���  �u �u�u�u�u�u�u�Ѓ�,]�U�졠��@H���  ]��������������U�졠��@H���  ]��������������U���u0�E�u,����u(�@H�u$��P  �u ���D$�E�$�u�u�Ѓ�,]����������������A    ����q�������@l�@��Y���������U�졠�V�@l��@�v�ЋM����u�A^]� �u����u�@lQ�u� ��3Ƀ������F^��]� �������������̋I��u3�á��Q�@l�@�Ѓ������U�������U��@lR�@�U�R�u�u�q�ЋM��U��;�u	�E���]� ���9U�D���]� �������U�졠��@H���   ]��������������U�졠��@H���  ]��������������U�������M�@�����   W��$�u���]��E�M�f/�w�Ef/�w(�����M�@���@,�$�u�Ћ�]����������U���0���W��M�Q�u�E��E��E��@�MЋ��   Q�M���~X�Ef/��~ �~P�Mv(��	f/�v(�f/�v(��	f/�v(�f/�wf/�v(��(ġ���E��U��]��@�M�@HQ�u�M�Ћ�]�������������U�졠��@H��0  ]�������������̋������������������������������̡���@H���  ��U�졠��@H���  ]��������������U���u0����u,�@H�u(���  �u$�u �u�u�u�u�u�uQ�Ѓ�0]�, ����U���u0����u,�@H�u(���  �u$�u �u�u�u�u�u�uQ�Ѓ�0]�, ���̡��Q�@H��,  �Ѓ�������������U�졠��u�@HQ��X  �Ѓ�]� �̡��Q�@H��\  �Ѓ�������������U��V�u��E�EP��������    ^]����������������U��QSV��MW�}3҉u��ϋ���t
����B��u��PSWV�M�)  �} ~(��   VW�}�W�M�  SVW�M��  _^[��]� ;�tSWV�M�l  _^[��]� ���U��V���v�������@l�@�Ѓ��Et	V���������^]� �����������U���V�u����   �ƙ+U��S��A�Z�W�	�<�ˉM��E��}�]���d$ �]��}�E���$    ��~I�����M��]��E��*�G���S����GN�C�u�}��W��~g�M��U����9u����    ���G���;�}��U;H}G���;�M��w������s��H�K�p�u�?��U;�~��M��N���_[^��]� ����̡��j �@Hh(  ���   Q�Ѓ������U��UV�u��+����� ~^�E�U]����S�ZW�]��I ��;�t7�]��$    �;H�}�p�ыH���H��H�P��p����;�u܋]�U�u���];�u�_[^]� ��U��QS�]W�}��+ǃ���M�=   ��   V�E��tu�7H�E��+����+����K��ǍǉU;�}9U|��;��;�}���9UL��M�PSW�u�   �u�M�S��V�u�z�����+������   �^_[��]� �M�SW�u�����^_[��]� ������������U��QS�]V�u;�t8W��F���;}$���N�M���
�H�@��J�R�;8|�E��:�B��;�u�_^[��]� U��ES�]VW�}�����9|���I ��;|�;�s$���p��O�H��w;�u����;�uǋ���_^[]� ���������̡��Q�@\�@�Ѓ���������������̡��Q�@\�@�Ѓ����������������U�졠��u�@\Q�@�Ѓ�]� �����U�졠��u�@\�u�@Q�Ѓ�]� ��U�졠��u�@\Q�@�Ѓ�]� ����̡��Q�@\�@�Ѓ����������������U�졠��u�@\Q�@ �Ѓ�]� �����U�졠��u�@\�u�@$Q�Ѓ�]� ��U���u����u�@\�u�@`�uQ�Ѓ�]� ������������U�졠��u�@\Q�@0�Ѓ�]� �����U�졠��u�@\Q�@@�Ѓ�]� �����U�졠��u�@\Q�@D�Ѓ�]� �����U�졠��u�@\Q�@H�Ѓ�]� ����̡��Q�@\�@4�Ѓ����������������U�졠��u�@\�u�@8Q�Ѓ�]� ��U�졠��u�@\Q�@<�Ѓ�]� �����U���SVW�}��j �ω]��������S�@\�@�Ѓ���S������3���~?��I ����M��@\Q�@`�MQh���V�u��Ѓ����u�U����u����K���F;�|�_^[��]� �������������U���S�]W�E��P���� ���}� |z���W�@\�@�Ѓ��E�P��� ���E���tWV3���~B�EP��� ���E�P��� ���M;M����Q�@\W�@�ЋMA���M;M�~�F;u�|�^_�   [��]� _�   [��]� ����������̡���@\� ������U�졠�V�@\�u�@�6�Ѓ��    ^]��������������̡��Q�@D�@$�Ѓ����������������U�졠�j �@D�u� �Ѓ�]��������U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�졠��@D� ]��U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�졠��u�@Dh2  � �Ѓ�]�����U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�졠�j �@D�u� �Ѓ�]��������U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�졠��u�@Dh'  � �Ѓ�]�����U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�졠��u�@DhO  � �Ѓ�]�����U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U�졠����@XQ� �M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ���������������U�졠����@XQ�@�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ��������������U�졠����@XQ�@�M�Q�ЋM�~ f��~@f�A�~@��f�A����]� ��������������U�졠���`�@XV�@WQ�M�Q�Ћ��E���   ���_^��]� �������������U�졠��u�@XQ�@�Ѓ�]� �����U�졠��u�@XQ�@�Ѓ�]� �����U�졠��u�@XQ�@�Ѓ�]� �����U�졠��u�@XQ�@�Ѓ�]� �����U�졠��u�@XQ�@$�Ѓ�]� �����U�졠��u�@XQ�@ �Ѓ�]� ����̡��j �@Dh�  � �Ѓ�����������U�졠�V�@@�u�@�6�Ѓ��    ^]��������������̡��Q�@D�@(�Ѓ���������������̡��Q�@D�@�Ѓ����������������U�졠��u�@D�u�@Q�Ѓ�]� �̡��j �@Dh:  � �Ѓ�����������U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U�������E�    �E�    ���   �U��@Rj�����#E���]�����������̡��j �@Dh�F � �Ѓ�����������U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U��E����u��]� �E�����E�    ���   �U��@Rj������؋�]� ̡��j �@Dh�_ � �Ѓ�����������U�졠�V�@@�u�@�6�Ѓ��    ^]���������������U��EV�0W�9;�t_3�^]� �P��u ��u9pu9qu��u�9yu�_�B^]� S�Y��u"��u9yu��u3��u/9pu*[_�   ^]� ��t��t;�u�P��t�A��t�;�t�[_3�^]� U���u�e������@]� ������������Vh��j\hD ����K  ����t�@\��tV�Ѓ���^�����U��Vh��j\hD ����K  ����t2�@\��t+V��h��jxhD �K  ����t�@x��t	V�u�Ѓ���^]� ���������U���Vh��j\hD ���fK  ����tG�@\��t@V�ЋEh��jdhD �E��E�    �E�    �0K  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh��j\hD ����J  ����t2�@\��t+V��h��jdhD ��J  ����t�@d��t	�uV�Ѓ���^]� ���������U��Vh��j\hD ���J  ����tZ�@\��tSV��h��jdhD �gJ  ����t�@d��t	�uV�Ѓ�h��jhhD �?J  ����t�@h��t	�uV�Ѓ���^]� �U��Vh��j\hD ���	J  ������   �@\��t{V��h��jdhD ��I  ����t�@d��t	�uV�Ѓ�h��jhhD �I  ����t�@h��t	�uV�Ѓ�h��jhhD �I  ����t�@h��t	�uV�Ѓ���^]� �����Vh��j`hD ���\I  ����t�@`��tV�Ѓ�^�������U��Vh��jdhD ���)I  ����t�@d��t	�uV�Ѓ�^]� �������������U��Vh��jhhD ����H  ����t�@h��t	�uV�Ѓ�^]� �������������Vh��jlhD ���H  ����t�@l��tV�Ѓ�^�������U��Vh��jphD ���yH  ����t�@p��t�uV�Ѓ�^]� ���^]� ���U��Vh��jxhD ���9H  ����t�@x��t	V�u�Ѓ���^]� �����������U��Vh��j|hD ����G  ����t�@|��tV�u�Ѓ�^]� 3�^]� ������U��Vh��j|hD ���G  ����t�@|��tV�u�Ѓ����@^]� �   ^]� ��������������U���Vh��jthD ���fG  ����tP�@t��tI�u�M�VQ�Ћu����P�`���h��j`hD �/G  ����th�H`��ta�E�P�у���^��]� h��j\hD ��F  �u����t4�@\��t-V��h��jdhD ��F  ����t�@d��th��V�Ѓ���^��]� �������U��Vh��h�   hD ���F  ����t���   ��t�uV�Ѓ�^]� 3�^]� U��Vh��h�   hD ���VF  ����t���   ��t�uV�Ѓ�^]� 3�^]� VW��3����$    �h��jphD �F  ����t�@p��t	VW�Ѓ������8 tF��_��^�������U��SV��3�W��    h��jphD �E  ����t�@p��t	VS�Ѓ������8 tph��jphD �E  ����t�@p��tV�u�Ѓ�������h��jphD �\E  ����t�@p��t	VS�Ѓ�����W���x�����tF�^����E_��t�0��~=h��jphD �E  ����t�@p��t	VS�Ѓ������8 u^�   []� ^3�[]� �����������U���Vh��h�   hD ���D  ����t<���   ��t2�u�M�VQ��h��j`hD �D  ����t�@`��t	�M�Q�Ѓ���^��]� �������U���Vh��h�   hD �ED  ����tS���   ��tI�u�M��uQ�Ћu����P�:���h��j`hD �	D  ����td�H`��t]�E�P�у���^��]�h��j\hD ��C  �u����t2�@\��t+V��h��jxhD �C  ����t�@x��t	V�u�Ѓ���^��]�������̋���������������h��jhD �oC  ����t	�@��t��3��������������U��V�u�> t+h��jhD �3C  ����t�@��tV�Ѓ��    ^]�������U��} W��t0h��jhD ��B  ����t�@��t�u�uW�Ѓ�_]� 3�_]� �������������U��Vh��jhD ���B  ����t�@��t�uV�Ѓ�^]� 3�^]� ������U��Vh��jhD ���iB  ����t�@��t�uV�Ѓ�^]� 3�^]� ������Vh��j hD ���,B  ����t�@ ��tV�Ѓ�^�3�^���Vh��j$hD ����A  ����t�@$��tV�Ѓ�^�3�^���U��Vh��j(hD ����A  ����t�@(��t�u�u�uV�Ѓ�^]� 3�^]� U��Vh��j,hD ���A  ����t�@,��t�u�uV�Ѓ�^]� 3�^]� ���U��Vh��j(hD ���IA  ����t�@0��t�u�u�uV�Ѓ�^]� 3�^]� Vh��j4hD ���A  ����t�@4��tV�Ѓ�^�3�^���U��Vh��j8hD ����@  ����t�@8��t�u�u�u�uV�Ѓ�^]� 3�^]� �������������U��Vh��j<hD ���@  ����t�@<��t	�uV�Ѓ�^]� �������������U��Vh��h�   hD ���F@  ����u^]� �u���   V�Ѓ�^]� ������U��Vh��h�   hD ���@  ����u^]� �u���   V�Ѓ�^]� ������U��Vh��h�   hD ����?  ����u^]� �u���   V�Ѓ�^]� ������U��Vh��h�   hD ���?  ����t�u���   �u�uV�Ѓ�^]� �����Vh��jDhD ���L?  ����t�@D��tV�Ѓ�^�3�^���U��Vh��jHhD ���?  ����t�u�@HV�Ѓ�^]� �U��Vh��jLhD ����>  ����u^]� �u�@LV�Ѓ�^]� ������������U��Vh��jPhD ���>  ����u^]� �u�@P�uV�Ѓ�^]� ���������U��Vh��h�   hD ���f>  ����u^]� �u���   �u�uV�Ѓ�^]� U��Vh��h�   hD ���&>  ����u^]� �u���   �u�u�u�uV�Ѓ�^]� ����������Vh��jThD ����=  ����u^Ë@TV�Ѓ�^���������U��Vh��jXhD ���=  ����t�u�@XV�Ѓ�^]� �U���Vh��h�   hD ���s=  ����tQ���   ��tG�u�M�Q���ЋuP���l���h��j`hD �;=  ����t|�H`��tu�E�P�у���^��]� h��j\hD �E�    �E�    �E�    ��<  �u����t3�@\��t,V��h��jdhD ��<  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh��h�   hD ���<  ����t���   ��t�u���u�u��^]� 3�^]� ������������U��Vh��h�   hD ���6<  ����t���   ��t�u����^]� 3�^]� ��U��Vh��h�   hD ����;  ����t���   ��t�u����^]� 3�^]� ��U��Vh��h�   hD ���;  ����t���   ��t�u����^]� 3�^]� ��Vh��h�   hD ���y;  ����t���   ��t��^��3�^����������������U��Vh��h�   hD ���6;  ����t���   ��t�u���u�u��^]� 3�^]� ������������U��Vh��h�   hD ����:  ����t���   ��t�u����^]� ���������U��Vh��h�   hD ���:  ����t���   ��t�u���u�u��^]� 3�^]� ������������Vh��h�   hD ���Y:  ����t���   ��t��^��3�^����������������U��h��jhD �:  ����t
�@��t]��3�]��������U���Vh��h�   hD ��9  ����u����u�HV�I�у���^��]Ë��   W�u�M�Q�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]���U��h���uhD �[9  ��]��������    �A    �A    �A    �����U��QV��~ uK���t����v�@<Q�@�Ѓ��    �~ t%�N��t������F�E��E�P�2������F    ^��]����U����E�VjP����������P�   �M���w�����^��]�U��EV��~ �Fu/h��jFj��������t�u��������3��F��u^]� �~ t3�9^��]� ����u�@<� �Ћȃ�3��ɉ�F   ��^]� ����V���F   ����@<�@��3Ʌ����^���������������U��	�����u	�@� ]� �@<�u�@Q�Ѓ�]� �����̃y t�   ËQ��u3�á��R�@<�1�@�Ѓ��������U��QV��~ uK���t����v�@<Q�@�Ѓ��    �~ t%�N��t�!����F�E��E�P�������F    ^��]����U��̴�����u�@� ]Ë@<�u�@Q�Ѓ�]�������U��̴��$V��u����A�0�����u�@<Q�@�Ћ�������I�E�ISP�ѡ���M�@Q�@V�С���M܋@Q�@�С��j �@j��@�M�h��Q�С���� �@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С������[t(�H�u�IV�ы���E�IP�I�у���^��]Ë@j�u��@H�M��С��j��@j��u�@L�u��M��С���u�@V�@�С��V�H�E�IP�ы���E�IP�I�у���^��]������������U��̴��$SV��u����A�0�����u�@<Q�@�Ћ�������I�E�IP�ѡ���M�@Q�@V�С���M܋@Q�@�С��j �@j��@�M�h��Q�С���� �@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С������t)�H�u�IV�ы���E�IP�I�у���^[��]Ë@j�u��@H�M��С��j��@j��u�@L�u��M��С���M܋@Q�@�С��j �@j��@�M�h��Q�С�����@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С�������?����@j�u��@H�M��С��j��@j��u�@L�u��M��С���u�@V�@�С��V�H�E�IP�ы���E�IP�I�у���^[��]���U��̴��$SV��u����A�0�����u�@<Q�@�Ћ�������I�E�IP�ѡ���M�@Q�@V�С���M܋@Q�@�С��j �@j��@�M�h��Q�С���� �@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С������t)�H�u�IV�ы���E�IP�I�у���^[��]Ë@j�u��@H�M��С��j��@j��u�@L�u��M��С���M܋@Q�@�С��j �@j��@�M�h��Q�С�����@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С�������?����@j�u��@H�M��С��j��@j��u�@L�u��M��С���M܋@Q�@�С��j �@j��@�M�h��Q�С�����@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С������������@j�u��@H�M��С��j��@j��u�@L�u��M��С���u�@V�@�С��V�H�E�IP�ы���E�IP�I�у���^[��]�����������U��̴��$SV��u����A�0�����u�@<Q�@�Ћ�������I�E�IP�ѡ���M�@Q�@V�С���M܋@Q�@�С��j �@j��@�M�h��Q�С���� �@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С������t)�H�u�IV�ы���E�IP�I�у���^[��]Ë@j�u��@H�M��С��j��@j��u�@L�u��M��С���M܋@Q�@�С��j �@j��@�M�h��Q�С�����@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С�������?����@j�u��@H�M��С��j��@j��u�@L�u��M��С���M܋@Q�@�С��j �@j��@�M�h��Q�С�����@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С������������@j�u��@H�M��С��j��@j��u�@L�u��M��С���M܋@Q�@�С��j �@j��@�M�h��Q�С�����@j �@@�M�Q�M�Q�M��Ѕ�����M܋@Q�@���С�����������@j�u��@H�M��С��j��@j��u�@L�u��M��С���u�@V�@�С��V�H�E�IP�ы���E�IP�I�у���^[��]���U��E�̴��EȉM]����������U�졠��@<�@]�����������������U��E����u��]�VP�M���(  �EP�E�P�M��E�    �E    �')  ����   �u�E���tA��t<��uX����u���   �@H�Ћ���ЋA���@xV���Ѕ�u+�   ^��]á���u���   �@T��VP�Y�������uՍEP�E�P�M��(  ��u�3�^��]��������U���DS3ۉ]�����M܋@V�@Q�С��S�@j��@�M�h��Q�С���M܋@<Q�@�Ћ�����I�E܋IP�у���u^3�[��]�WV�M�3���'  �E�P�E�P�M��	(  ���  ��}���   ����u����   �@T�Ћ�������   ������A�M̋@Q�С�����@�M̋��   Qj�M�Q���Ћ�����I�E܋IP�ы���A�M܋@QV�С���M��@Q�@�С�����@�u�@x�M����E���t�E� ��t����M܋@Q�@����Ѓ���t����M̋@Q�@����Ѓ��}� u!�E�P�E�P�M���&  ���������_^[��]Ë}���_^[��]��������������U���@SV�u3ۉ]���u^����M��@Q�@�С��V�@j��@�M�h��Q�С���M��@<Q�@�Ћ�����I�E��IP�у���u^3�[��]�V�M��&  �E�P�E�P�M��E&  ��t�W�}�E�����   ����u����   �@T�Ћ�������   ������A�MЋ@Q�С�����@�MЋ��   Qj�M�Q���Ћ�����I�E��IP�ы���A�M��@QV�С���M��@Q�@�С�����@W�@x�M����E��t�E ��t����M��@Q�@����Ѓ���t����MЋ@Q�@����Ѓ��} tA�E�_^[��]Ã�u2�M���t+���Q���   �@H�Ћ���ЋA���@xW���Ѕ�t��E�P�E�P�M���$  �������_^[��]�������̡���@<�@�����U��Q�=Դ uX�̴��t!����5ܴ�@<Q�@�Ѓ��̴    �ش��t#蹹���ش�E��E�P�(������ش    ��]���������t������������t�����������U��QV���t�j ��E�P�u��ӵ����^��]�����������̡���@��  �ࡠ��@��(  ��U�졠����@�U䋀   R�ЋMP轸���M�������E��]� �����������̡���@��$  ��U�졠��@��  ]��������������U�졠��@���  ]�������������̡���@��  ��U�졠��@���  ]��������������U�졠��@��x  ]��������������U�졠��@��|  ]�������������̡���@��d  ��U�졠��@��p  ]��������������U�졠��@��t  ]��������������U���EV���t�t	V��������^]� �������������̡���@��   ��U�졠�V�@�u��$  �6�Ѓ��    ^]������������U�졠�V�@��(  V�u�Ѓ���^]� ������������U�졠�Q�@�u��,  �Ѓ�]� ��U�졠�Q�@�u��,  �Ѓ����@]� �������������U��E��t�P�3ҡ��R�@Q��8  �Ѓ�]� ������U�졠��u�@Q��<  �Ѓ�]� ��U���u����u�@�u��@  Q�Ѓ�]� ������������U�졠��u�@�u��D  Q�Ѓ�]� ���������������U�졠��u�@Q��H  �Ѓ�]� ��U�졠����@V��L  W�uQ�M�Q�Ћ���}�IW�I���ы��W�IV�I�ы���E��IP�I�у���_^��]� ������������̡��Q�@��T  �Ѓ������������̡��Q�@��P  �Ѓ�������������U�졠��u�@Q��X  �Ѓ�]� ��U�졠��u�@Q��l  �Ѓ�]� �̡���@��0  �ࡠ��@��4  �ࡠ��@��p  �ࡠ��@��t  �ࡠ��@��\  ��U�졠�V�@�u��`  �6�Ѓ��    ^]������������U���u����u�@�u��d  �u�uQ�Ѓ�]� ������U���u����u�@�u��h  �u�uQ�Ѓ�]� �����̡��Q�@�@�Ѓ����������������U���u����u�@�u�@X�uQ�Ѓ�]� ������������U�졠��u�@Q�@\�Ѓ�]� ����̡��Q�@�@ ��Y�U�졠����@V���   h�  Q�M�Q�Ћ��P���   �@8�Ћ�������   �E��	P�у���^��]��������������U�졠��@��   ]��������������U���u����u�@�u�@Q�Ѓ�]� ���������������U���u����u�@�u���   �uQ�Ѓ�]� ���������U�졠��@�@$]�����������������U���u����u�@�u�@(�uQ�Ѓ�]� ������������U���u����u�@�u�@,�uQ�Ѓ�]� ������������U���u(����u$�@�u �@`�u�u�u�u�u�uQ�Ѓ�(]�$ �������������U�졠�V�@W�@��W�Ћ��W�J���I���u����u�Q�u�N�QHP�B4j j W�Ѓ�(_^]� ���������������U���u ����u�@�u�@4�u�u�u�uQ�Ѓ� ]� ���U�졠��u�@�u�@@Q�Ѓ�]� ��U�졠��u�@Q�@D�Ѓ�]� ����̡��Q�@�@L�Ѓ���������������̡��Q�@�@L�Ѓ���������������̡��Q�@�@P�Ѓ����������������U�졠��u�@Q�@T�Ѓ�]� �����U�졠��u�@Q�@T�Ѓ�]� ����̡��Q�@�@h�Ѓ����������������U�졠��u�@�u���   Q�Ѓ�]� ���������������U�졠����@V�u���   �uQ�M�Q�Ћuj �    �F    ���P���   V�I�ы���E����   P�	�у� ��^��]� ��������̡���@� ������U�졠�V�@�u�@�6�Ѓ��    ^]���������������U���u����u�@�u���   �u�uQ�Ѓ�]� ������U�졠�V�@�u�@�6�Ѓ��    ^]���������������U��QS�]V�C    �����@V�@h�Ѓ���u9h�h  hx�h  @谀�����=�� t
�=�� t�^3�[��]� ����M�Q�MQ�u�E    �@V���   �Ѓ���t�3�9u�~%W�E�<� �<�tj���)  ��t��F;u�|�_�E�E�EP�������   ^[��]� �����������U��QS�]V�C    �����@V�@h�Ѓ���u9h�h)  hx�h  @�������=�� t
�=�� t�^3�[��]� ����M�Q�MQ�u�E    �@V���   �Ѓ���t̃} t�3�9u�~<W�E����t*���Q�@�@h�Ѓ���t�Ej�<����*  ��t�8F;u�|�_�E�E�EP�������   ^[��]� ��������������U�졠��@��x  ]�������������̡���@��|  ��U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]��������������U�졠��@���  ]�������������̡��Q�@���   �Ѓ�������������U�졠��u�@Q���   �Ѓ�]� �̡���@���   ��U�졠�V�@�u���   �6�Ѓ��    ^]������������VW���O�Ī��W�f�G f�G(f�G0f�G8f�G@f�GHf�GPf�GX�    �G`    �Gd    �Gh    �Gp�Gx�����G|   ��_^�������V���X   �N^�?������������������W��    �A`    �Ad    �Ah    �Ap�Ax�����A|   ���������������SW�����t7�������xP t$V������j j �pPj�GP���}����H ���^�    �O`��t���Q�@�@�Ѓ��G`    _[��������������h�h�   h�   謦������t������3�������������U��S�]W�;��tV�7�u��t6��������xP t#��������Mj j �pPj�GP������H ����    �O`^��t���Q�@�@�Ѓ��G`    �O�ک����E�EP�L������    _[]����������������U�졠�S�@V��   W��W�_dS�wx�w`�uV�Ѓ��G|����   �? ��   �; ��   �wpV�_hS�u��_������u8h�h)  W�hx�h  @����z�����=�� t
�=�� t��u�O辬�����������xP u����"������j j �pPj�GP�������H ��ЉG|��t��������G|_^[]� �G|�Gx����_^[]� �G|�����    ����6�@�@�Ѓ��    �G|_^[]� ���������������V���x���W��    �F`    �Fd    �Fh    �Fp�Fx�����F|   ^������U��QW���d �G`t~S�];_xttV�7�ΉE�u�������xP u����#�������M�S�u�pPj�GP�����H ��ЉG|^��u�E�_x��t�    �G`[_��]� �M�Gx������t�3�[_��]� �����������U��E��t	�Ap� �yd t�Ah]� 3��y|��]� ���U���u ����u�@�u�@�u�u�u�uQ�Ѓ� ]� ���U�졠��u�@Q�@�Ѓ�]� ����̡��Q�@�@��Y�U�졠��u�@�u�@Q�Ѓ�]� �̡���@� ������U�졠�V�@�u�@�6�Ѓ��    ^]���������������U��VW���T����u���u�x@�u�A����H ���_^]� ����U��VW���$����u���u�xD�u�����H ���_^]� ����W��������xH u3�_�V��������ύpH������H �^_�����U��W��������xL u3�_]� V�������u���u�pL�u�����H ���^_]� U��W�������xP u���_]� V���o����u���u�pP�u�u�Y����H ���^_]� ������������U��W���5����xT u���_]� V�������u���u�pT�����H ���^_]� ��U��W��������xX u���_]� V��������u�ύpX������H ���^_]� �����U���SVW�}�م�t.�M�������������pL�E�P�������H ��ЍM�� ����u��tW����M��@Q�@�С���M��@V�@Q�С���M��@Q�@�Ѓ����;����H@��t���V�@Q�@�Ѓ�_^[��]� ���������U��VW�������u�΍xH������H ���_^]� ����������U��W��������x` u
� }  _]� V�������u�ύp`�����H ���^_]� ���U��SVW�������x` u� }  �#�������p`�E���P���l����H ��Ћ�����]�IS�I�у�;�>���S�@�@�Ѓ�;�)���.����u���u�pDS�u�����H ���_^[]� _^�����[]� U��W��������xP u
�����_]� V��������u���u�pP�u�u�u�u������H ���^_]� ����U��W�������xT u
�����_]� V�������u���u�pT�}����H ���^_]� U��W���e����xX tV���W����u�ύpX�J����H ���^_]� �������������U�졠���   �@V� ���Љ���3  S�u�M��¡������M��@Q�@�С��j �@j��@�M�hP�Q�Ѓ��E�P�M�舡���E�P�E�P��d���P�t�����P�E�P�ǥ����P�E�P躥�����j �ЋAj��@R�6�Ѓ����M���財���M�誡����d���蟡���M�藡������M��@Q�@�Ѓ��M��{��������[t�@�6�@�Ѓ��    ��^��]� �E�M�Q�E�   �E��@jd�6���   �С���M����   Q� �Ѓ���^��]� ��U���V�E�P�u���E�    �E�    �E�    �E�    �E�    �E�    �A4  ����t�}� t�M��\o�����^��]� �    ��^��]� �̡��V�@��@�6�Ѓ��    ^����U����E�P�u�E�    �E�    �E�    �E�    �E�    �E�    �3  ����t*�}� t$�E�~E�f� �~E�f�@�~E�f�@��]ËE�     �@    �@    �@    �@    �@    ��]����U����E�P�u�E�    �E�    �E�    �E�    �E�    �E�    �3  ����t�}� t�M��/n����]�3���]������U��USV��W�F��~���;�~W��@�+����ׁ�  �yJ���Bu��u	�   +��hX�h  ��    PQ耛���Ѓ���t�N��~��_�^^[]� �F_�F^��[]� ��̸   � ��������3�� �����������3�� ����������̸   @� ��������3�� ����������̸   � ��������U�졠��u�H�I�ыE��]� ��̸   � ��������U����   V�u��u3�^��]�h�   ��@���j P��O  �E�E��E�E��Eh�   ��@�����@���P�u��`����uǅD���бj�E����E����E����E����E����E����E����E����S���� ^��]��������U����   h�   ��@���j P�$O  �Eh�   �E���@���P�uǅ`���    �uj��R���� ��]�����U���   SV�u(W3�3��]����w  ����M�@�@<�Ѕ��F  �5����E�����   �EP�M�莜������M�@Q�@�С��W�@j��@�M�hP�Q�Ѓ��E�P�M��U����u�Wj��E�P�E�P��\���P�_?�8�����P��x���P舠����P�E�P�{�������P�P����E���t�E� �� t�M�����s�����t��x�������`�����t��\�������M�����t�M̃���=�����t����M�@Q�@����Ѓ���t�M������}� t�u(�u$�u��u�u�u���������E�P�	������V�u$j �u�u�u�p�����������E�IP�I�у���_^[��]Ë�`��`��`��`��`��`��` ��`�����U��EH������   �$����   ��]á��@�������   �u��l����=�:  }	�������]Ã} t�E�Pj�E����E�o   �E�    ��S������t{���
�������tu�u��藞���   ��]��u�u�C����������H��]�������]����u7������������t#蚚�����E�EP�	�������    �   ��]Ã����]���|�������b�����U���Mu�E���E���   ]� ���������������U��� �@�V���.�vf(�fT �f/�f(�fT ��U��M��M��%  f/��  ���f/�vFf/�v@�,��,���   ��$    ������ʅ�u�fn�����^��^��.�v^��]�f/�v(��(����^��%��f/�v1(��Y��Y��Y��E�(��Y��.�v(��M��M�f/�v(��E��E��f��    �E��E���i  �]��E�f/(��M��M��E��E�s���^���F�^��F^��]�W������F^��]��������U���E� �f/�V��w��f/�v(��Y�����X(��E�E�$�#c  ���������F�
�����^]� ���U����M�U3�W�f/�fT ��X(���3�f/�V����3��M��E�;������$�M�b  ��EfT ��E�X(��E�E�$�b  ����]�E��f/��Fv9h��j!hx�h  @�i�����=�� t
�=�� t�����F�} u�fW0����������^��]� ��U���E���f/�V���Fv9h��j/hx�h  @�h�����=�� t
�=�� t�����F^]� ����U���M�����f/�V��v9h��j8hx�h  @�.h�����=�� t
�=�� t�����M��Y����E��E��$�0a  �]��F�$�"a  �E��]��^E��E��E��$�a  ��E�$��`  ���^�������^��]� ����U�졠�Q���   �@X�Ћȃ���u]� ����u�@|�u�@Q�Ѓ�]� ����U�졠�Q���   �@X�Ћȃ���u]� ����u�@|�u�@8Q�Ѓ�]� ����U��UV��j ����j �@j �@R�Ѓ��F��^]� ���̡��V�@j �@j ��j �6�Ѓ��F^�U��V��N��u3�^]� ���Q�u�@�u�@�6�Ѓ��F�   ^]� ������U��M�]�`����U��M�]�`����V��h���d��F    ���V�@Ph`�� hP��Ѓ��F��^����������̃y �d�u����q�@P�@��Y���U��I��u3�]� ���j �u�@P�u�@Q�Ѓ�]� ���U��I��t����u�@PQ�@�Ѓ�]� ��������������U��I��t����u�@PQ�@�Ѓ�]� ���������������    �A    ���V����t&���Q�@P�@L�С���6�@P�@<�Ѓ��    ^����������������U��SVW�����t���Q�@P�@<�Ѓ��    �G    �M�]h��S�O���h`��@PhP��@8Q�u��3����9u~E���x u�@   ����HP���p�A�Ѓ����V�@P�7�@@�Ћ�F���A;u|�3�9_^��[]� �����������U���u�E�u�p�,���]� ��������U��SVW��3�9w~=�]���V�@P�7�@@�ЋЃ���t-���j �APS�@jR�Ѓ���tF;w|�_^�   []� ����7�@P�@L�Ѓ�3�_^[]� ������������̡���1�@P�@D�Ѓ��������������̡���1�@P�@H��Y���������������̡���1�@P�@L��Y���������������̡���@P�@P�����U�졠��@P�@T]����������������̡���@P���   ��U�졠��@P���   ]��������������U��M�]�`����U��V��~ �d�u����v�@P�@�Ѓ��Et	V�_�������^]� �����3���������������U��M�EQ��Ej�u�A�tP����]���������������̸   �����������U��V�u��t���u6j�u�uP������u3�^]Ë���O���ȅ�t��t��E3�;AOʋ�^]�������U��j�u�3P������u]Ë��O�������]�������������    �A    �A    �A    �����U��QV���E��E�P蛌���    �F�E��E�P膌���F    ���F    �F    ^��]����������U��V��W�}�    �F    �F    �F    �Gj;Gu2j�   ��tY�����G�A��G�A�F_�    ��^]� j�   ��t'�����G�A��G�A��G�A�F�    _��^]� �����U��V�u���    �F    �F    �F    �  ��^]� U��V�u���r  ��^]� �����������U��QSV���E��E�P�Z����    �F�E��E�P�E����]���F    �F    �F    ����   �ÙW�ȋ��������;�u;�uh��jIQ車�����3����tV�}��tZ�Ǚ�ȋ������E���;�u9Uuh��jNQ�}������3��F��u"��E�EP衊�����    _^3�[��]� �~_�^^�   [��]� ^3�[��]� ���������������U��QV���E��E�P�K����    �F�E��E�P�6����F    ���F    �F    ^��]����������U���V��W��E��E�P������    �F�E��E�P�����}���F    �F    �F    ����   �? ��   �G����   �S�ȋ��������;�u;�uh��jlQ�'������3��[��tF� tJ�G��tC����M�Q��RP�E���E�q   �E�    �������F��u�������_3�^��]� �G�F�G�F��P�7�6��7  �N����t�F��P�wQ�7  ��_�   ^��]� ������U���SV��W��E��E�P�ǈ���    �F�E��E�P貈�����} �F    �F    �F    �  �}���  �Ǚ�ȋ��������;�u;�uh��h�   Q��������3����tG�]��tS�E��tL����M�Q��RP�E���E�   �E�    ��������F��u������_^3�[��]� �E�F�3�E�Pj j�F   �E���E��   �E�    �������F��t���    P�u�~�6�m6  ����t!�F��PS�v�V6  ���   _^[��]� �F�8_^�   [��]� ���    �A    �A    �A    �����U������   �U��V�HWW�3��<��D$�|$@�L$}
��_^��]� ����  �0�U�f(ύ@�F�~ʍ@f(��D��,��t��\D��D$�\t��8�L$(�|$ �T$�\$0�\��D$8����   ��������f(ƍ@f(��$��T��\T��\��\��\\����Y��Y��Y��Y��\�f(��Y��Y��XL$(�\�f��\$0�\��L$(�Xl$�Xt$ �l$f�f(��D$ f�O�f����T$W��(��YL$(�YD$ �}f�?�X�f(��Y�f�f��X��`Z  �T$(�\$ f(�W�f.͟��Dz�L$f(�f(�f(��&����^��L$f(�f(��Y��Y��Y�f�gH�% �fT�fT�f/�f�wPf�GX��   f(�fT�f/���   �GH�WX�gP(��Y�(��Y��\��Y��\�f�_�\�f�O f�g(�OX�P�Y(�W�gH(��YG (��YWP�\�(��YG(�Yg �Y�f�0�\��\�f�_8f�g@�)  �WPfT�f/��_X��   �OH�Y�f(��Y��\��\��Y�f�Gf�_ �\�f�O(�(�G �YGX�YP�O�wH(��Y_X�YOP�\�f(��YG(�Yw f�0�\��\�f�_8f�w@�   f(��Y�(��Y��\��GH�Y�f�O0�\��\�f�_8f�G@�oP�X�Y8�OH�w0(��YG@(��Y_@�YO8�\�(��YGX�Y�f��\��\�f�_ f�w(�D$`WP��  �U���D$�   ���W�3�3Ʌ�~w��r]�p��W�W�%  �yH���@��+���    �o���f���oD��f��;�|�f��fo�fs�f��fo�fs�f��f~ϋt$;�}�F<�A;�|���t$�M��u�A0�D$(���q �@�D$    ���d��\��Y�f(��YI�D$(�Y��X	�D��Xq�@�X��AH�Y��X��A8�Y��L$ �I(�X��AP�Y��Y��T��X��A@�XI�Y��$��X��AX�Y�(��YY�X�(��YA0�Xf�L$X�L��D$�X�(��YAH�@���X�(��YA8�YQ@�\$(��YY �Ya(�D$�XY�Xa�X�(��YAP�YIX�X��X��X��\$0f�d$8���  3�������|$�D$(׋��@�,��T��L�f(��Ya(��YA0�X!f(��YY �Yi(�X��XY(��YAH�Xi�D$@�X�(��YA8�YQ@�D$�X�(��YAP�YIX�X��T$0�X��X�(�f(��\��\��\�f�\$0�YD$�YL$ �Y��X��~D$�D$ �~D$8f�D$X�X�f�f�d$f�l$8�X�;D$������|$@�D$@_^��]� ������������U�������������U�   @t������@��wg�$���E� ����E� ���]� �
�E��E�J�]� �J�E��E�J�]� �J�E��E�J�]� �J�E��E�
�]� ����������������U��S��V�����%���W��   @t�����ʃ��};�t�����t�u�����t��u;�t?�����t7�΁����Eǃ��t����   �_�^�[]� ��   ���Ё�   @�_^[]� �U�������AW�SVf(�f(�f(�W�L$�\$�T$ �D$���L  �9�u������Ш�)  ���������U��Z�@�[�<��l��\<��\l�;Zuc�\��B�\\��@�d��\d��T��\T��4��\4�f(��Y�f(��Y��Y��\�f(��Y��\��Xd$(��d�d��B�\d��@�B�@�T��\��\\��\T��4��\4�f(�f(��Y��Y��Y��\�f(��Y��\��X\$�XL$�Y��Y��\$�L$�\��Xt$ (��T$ ���L$�����f(��Y�f(��Y��X�f(��Y��X��R  f(�W�f.П��D�Ez� �@�@_^[��]� ����^�_^[(��YD$� (��YD$�@�D$�Y��@��]� ���������U���<����5���A3�f�f�f�f��E��M��}��u��m��e�U�E����  S�V�uW�������Ш�v  ���������M��@��tn��f/�v	f(��E��\�f/�v	f(��M��\�f/�v	f(��}�f/�v	f(��u��T�f/�v	f(��m�f/�vIf(��>�~4��~l��~d�f�f�f�   �u��m��E��M��}ԉU��e�A�@��tn��f/�v	f(��E��\�f/�v	f(��M��\�f/�v	f(��}�f/�v	f(��u��T�f/�v	f(��m�f/�vIf(��>�~4��~l��~d�f�f�f�   �u��m��E��M��}ԉU��e�y���tn��f/�v	f(��E��\�f/�v	f(��M��\�f/�v	f(��}�f/�v	f(��u��T�f/�v	f(��m�f/�vIf(��>�~4��~l��~d�f�f�f�   �u��m��E��M��}ԉU��e�A;�t0�@�Mč�P�  �U��e��m��u��}��M��Eă��M��m���_^[��tb�Ef(��X�f(��X��(�f(��X��Y��Y��Y�f�f�Pf�H�\0�\h�\`�Ef�0f�hf�`��]� �EW�f� f�@f�@�Ef� f�@f�@��]� ��������̋Q3���|�	��t��~�    t@��Ju��3�����������U��QV�u��;�}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}���x(���t"�v3Ʌ�~�I ���%���;�tA��;�|�_���^]� _��^]� ���������U��SV�q2ۅ�~:�W�}�
����%���;�u��   @u�����t	�   ���3�
؃�Nu�_��^��[]� �������������V�q3҅�~�	�d$ ��   @u	�����tB��Nu��^�����V�q3҅�~�	�d$ ����ШtB��Nu��^�����������U���V��3�9N~�A�d�����;N|��N��~jS�   3�W�U��]�����x9���������;�}*������<����������;�u��   ��@;F|ۋU��]��NB���B��]��U�;�|�_[^��]�����������h��jh_� ���������uË@����U��V�u�> t/h��jh_� ��������t��M�@�MQ�Ѓ��    ^]���U��Vh��jh_� ���y�������t�@��t�u����^]� 3�^]� ��������U��Vh��jh_� ���9�������t�@��t�u����^]� 3�^]� ��������U��Vh��jh_� �����������t�@��t�u���u�u��^]� 3�^]� ��U��Vh��jh_� ����������t�@��t�u����^]� 3�^]� ��������U��Vh��j h_� ���y�������t�@ ��t�u����^]� 3�^]� ��������U��Vh��j$h_� ���9�������t�@$��t�u����^]� 2�^]� ��������Vh��j(h_� �����������t�@(��t��^��3�^������Vh��j,h_� �����������t�@,��t��^��3�^������U��Vh��j0h_� ����������t�@0��t�u����^]� 3�^]� ��������U��Vh��j4h_� ���Y�������t�@4��t�u���u��^]� ���^]� ����Vh��j8h_� ����������t�@8��t��^��3�^������U��Vh��j<h_� �����������t�@<��t�u����^]� ���������������U��Vh��j@h_� ����������t�@@��t�u����^]� ���������������U��Vh��jDh_� ���i�������t�@D��t�u����^]� 3�^]� ��������U��Vh��jHh_� ���)�������t�@H��t�u����^]� ���������������Vh��jLh_� �����������t�@L��t��^��3�^������Vh��jPh_� ����������t�@P��t��^��3�^������Vh��jTh_� ����������t�@T��t��^��^��������Vh��jXh_� ���\�������t�@X��t��^��^��������Vh��j\h_� ���,�������t�@\��t��^��^��������U��Vh��j`h_� �����������t�@`��t�u���u��^]� 3�^]� �����U��Vh��jdh_� ����������t�@d��t�u���u��^]� 3�^]� �����U��Vh��jhh_� ���y�������t�@h��t�u���u�u�u�u��^]� ���U��Vh��jlh_� ���9�������t�@l��t�u���u�u��^]� 3�^]� ��U��Vh��jph_� �����������t�@p��t�u���u��^]� 3�^]� �����U��Vh��jth_� ����������t�@t��t�u���u��^]� 3�^]� �����U��Vh��jxh_� ���y�������t�@x��t�u���u��^]� 3�^]� �����U��Vh��j|h_� ���9�������t�@|��t�u����^]� 3�^]� ��������U��Vh��h�   h_� �����������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh��h�   h_� ����������t%���   ��t�u���u�u�u�u�u��^]� ���^]� ��U��Vh��h�   h_� ���V�������t%���   ��t�u���u�u�u�u�u��^]� ���^]� ��U��Vh��h�   h_� ����������t���   ��t�u���u�u�u��^]� 3�^]� ���������U��Vh��h�   h_� ����������t���   ��t�u����^]� 3�^]� ��U��Vh��h�   h_� ���v�������t���   ��t�u����^]� ���������U��Vh��h�   h_� ���6�������t���   ��t�u���u��^]� 3�^]� ���������������U��Vh��h�   h_� �����������t���   ��t�u���u�u��^]� 3�^]� ������������U����M�U�E�R�X�A�\B�\��\Y�Y �Y�Y�X��X��U��E���]�����U��h���uh_� �K�����]�������U����   �M�qX�I8�y(�A@�YAP�Y�f(��YQP�E��M��\��A �E��Y�f(��U��Q �YQ@�\��E�(��YA8�U��M��}��E�(��Q0�\��A�Y��Y�W��]��e��X��AH�Y��X����f.џ��DzB�Ef�f�@f�H0f�HHf�Hf�H f�@8f�HPf�Hf�H(f�H@f�@X��]��^��y�E��A(��Y�(��Yq@(��Ya8�(��YYP(��Yy �\��e�(��\��e��YA0�\e��YIH�\u��\��i�X��E��\E��Y��Y��Y��Y�V�X�W�YM���8����I�YM�(��\��\��YAH�Yy0�X��X��]��Y���@����E��\E��Y��QH(��YI@�X��E��Y��X��y0��P����E��Y��Y���X����E��Y���H�����`���(��YAX�\�(��YA(�Y���h���(��YIX�\��Y���p���(��YA@(��YI(�E��8������\�(��YA8�YU��Y���x���(��YIP�Y}��\�(��Yi8�YAP�Y��\��\й   �M��Y��Y��m��U��_^��]��U��y0 �Etr��f/�v�	�H�Af/�v�I�H�Af/�v�I� f/Av�A�@f/A v�A �@f/A(vJ�A(]� �~ f�A�~@f�A �~@f�A(�~Af��~A f�A�~A(f�A�A0   ]� �������������U��h�jh�f �L�������t
�@��t]�����]�������U��Vh�jh�f ����������t=�~ t7�u8�E�u4�u0�u,�u(����P�l���u�F�Ѓ�4�M���l����^]ÍM����l����^]������U��h�jh�f ��������t
�@��t]��3�]��������U��h�jh�f �|�������t
�@��t]��3�]��������U��h��uh�f �K�����]�U��V�u���W.  �����^]� U��V�u���<.  �����^]� U��V�u���!.  �����^]� U��V�u���.  �����^]� ����.  �.  U��V�������-  �EtV��#��Y��^]� U��V����-  �EtV��#��Y��^]� U���j�E�P�M��E����o-  h p�E�P�E���b.  �U����E�E�EP�M��-  htp�E�P�E����4.  �U����E�E�EP�M���,  h�p�E�P�E����.  �U��=4� �0�t�M9t���x u�3�]Ë@]�U��=�� ���t�M9t���x u�3�]Ë@]�WhT���� ���uV�(�V��  ��Y����|�^��_�U��EV����u	j�X=  ���}k�(�P�  Y��^]� hT��$���yV�(�V�g  ��Y����|�^Ë��u	j�i>  YÃ�}k�(�P�j  Y��IG  U��V��N  �ujh   ���T  YY�F��th   ��K  P�v��  ���F   ��K  �f �F�N  �@�F��t
P�*N  Y�F��^]�U���V�uW��u�N  �x�XN  ��~��E���u�E�H�����   �� �   S�]��   s��uS�rM  Y��u�   �F�Xtx��u�����E��K  �U����H% �  ��F�������H������tj�U�]�E X�
3��]�E @j�u��M�jQP�EPh   Wj �hS  ��$��u������E�t	�M����[_^��U���V�uW��u�M  �x�[M  ��~��E���u�E�H�����   �� �   S�]��   s��uS�L  Y��u�   �F�Xtx��u�����E��J  �U����H% �  ��F�������H������tj�U�]�E X�
3��]�E @j�u��M�jQP�EPh   Wj �kR  ��$��u������E�t	�M����[_^��U��EV��3ҍN�F   �4�V�V�V�Fh@��Q�k   ��^]� �I��P��t�j����V���Σ�������V�r��Y�5����u�^�V��V�4�9  �~ Yt	�v�&  Y�f �P�^�U��SW�}��9;t>�; t�3�&  Y�# ��t*�? V��tF�> u�+�FV��0  Y���tVWP�  ��^_��[]� U��V���v����EtV����Y��^]� U��j���Y��t�����M�H�3����]á���j����8  j �M������5���e� ��u;V�  ��V�'  YYhD�N�F?   �����5������P�������} t����P�M��������I8  �j���P8  j �M��A����}�e� �w��GN����t��P��t�j�����u��w�?%  Y�M��`�����7  �U��j j �Q  YY��u���V�uP�N$�f����} t�uj �qQ  YY��u�@P�N,�B���^]�U��E�x$ t�p$j �DQ  YY]�U��j �5��Y��t�u���k���]�3�]�U��=�� uh�����|  Y�E���]�U��E���t��P��t�j���]�U��Qj �M��%���h��������%�� Y�M��g�����U��Qj�M�������M�A   �Q������t;�t�B�A��r�A�����A�M����������U��VW���w,��vW�u�V�6����u�_^]� U��V�u�F��t�����������   �v0��t�����V���Y^]�VWj �������G(��t�0P���Y�ƅ�u�G,�g( ��t�0P����Y�ƅ�u�g, _^�U��EVW3ɋ��Ѓ���   A�@t��t��%;���3�;�t���F��u��<�� u3��T��t!�
t�uj �u�L   ����t	P�;  Y���uV�u�0   ������t�tjj V�SR  ����tV�ˋ�_^]�U��]�U���U���u�E�4�P�u��P  ��]�U���u�0�]�U��j h�  �u��R  ��]�U���u�(�]�U���u�,�]�����AP����<���t�Ћ����
r��U�졀�����U  �uH����8�������]��5���<���t��j���  jj �6U  ���MU  Vjj ��L  YY��V�8���������ujX^Ã& 3�^�jhq��  蓊  �e� �u�#   Y���u��E������   ���/�  Ëu��n�  �U��QSV�5<�W�5�����5���E��֋؋E�;���   ��+��O��rvP�f�  ���GY;�sG�   ;�s�Ƌ]��;�rPS��L  YY��u�F;�r>PS�L  YY��t1��P���8�����u�8��KQ��8�����E�3�_^[��U���u����������YH]�U��V�u��t�U��t	�M��u��OU  j^�0�;�  ��^]�W��+���A��tJu�_��u��"U  j"��3���WV�t$�L$�|$�����;�v;��h  �%Ⱦs��  ���   ��  ��3Ʃ   u�%���  �%Ⱦ ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf����8����   u������r*��$�8��Ǻ   ��r����$�L�$�H��$���\��#ъ��F�G�F���G������r���$�8�I #ъ��F���G������r���$�8�#ъ���������r���$�8�I /����D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�8��HP\p�D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$�������$���I �Ǻ   ��r��+��$���$����4�F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I ���������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��������D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̋L$�D$WSV�=ľ��  ��   ��������   fn��p� �f�����������t��   u�foft�f�څ�u�   f~ڻ�  #؁��  w'�of��ft�ft�f��f�ك���t��ۃ�����tj��:�u��ЍN��  ��u9#ځ��  w/�o
foft�ft�ft�f��f�څ�u�������������t:�b��������H^[_�3�^[_À9 t�����  #ف��  w�o�"�   �1��f: �fs�Kt	��t����f~»�  #؁��  v���t�:�t�����f:c@�w�s�����׋��  #ށ��  w)��  #ځ��  w�o
����f:cN�q�y��L�������A���:�x�������뭊����to�q��tU���L$���:�t��t���:�t
��u�^[_3�Ê��:�u�~��a��t(���:�u��A��t�f���:�t��3�^[_���X�  �G�^[_Ë�^[_�U��V��M�F ��uf�ɓ  �ЉV�Jl��Jh�N�;��t����Bpu�i�  ��F; �t�N����Apu�̍  �F�N�Ap�u���Ap�F�
���A�F��^]� U��QQ�H�3ŉE�SV�u��u��K  j^�0讄  �3  �uV�K�  YY;Er� �׋U����   ��tJj�p3�SSj�Vh   QR�A  �ȃ�$�M���u2�fK  � *   �[K  � ��   �<a|<z, �F�> u�3��   9Ms��-K  j"�f�����~Ej�3�X���r9����   w���J�  �܅�t���  �Q�X   ��Y��t	���  ���M���u��J  �    �i����Uj��pQSj�Vh   ���   R�@  ��$��tS�uV�)��������
�J  j*^�0S�   Y�ƍe�^[�M�3���   ��U��E��t���8��  uP�d  Y]�U��=� u;�E��u�7J  �    �"�  3�]À8 ��t+���a|
��z�� �A�9 u�]�j j��u�   �E��]�U��j �u�u�   ��]�U����u�M��g����E�P�u�u��������}� t�M��ap���;H�u����  ����WV�t$�L$�|$�����;�v;��h  �%Ⱦs��  ���   ��  ��3Ʃ   u�%���  �%Ⱦ ��  ��   ��  ��   ��  ��s����v����s�~���vf����   tc����   foN�v�fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�   foN��v��I fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v�VfoN��v���fo^��0foF fon0�v0��0fo�f:�ffo�f:�fGfo�f:�fo �0}��v��|�o���vf�����s����v����s�~���vf���������   u������r*��$����Ǻ   ��r����$���$����$�L��,#ъ��F�G�F���G������r���$���I #ъ��F���G������r���$���#ъ���������r���$���I �����|tl�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���������D$^_Ð���D$^_Ð���F�G�D$^_ÍI ���F�G�F�G�D$^_Ð�t1��|9���   u$������r����$�T�����$��I �Ǻ   ��r��+��$�X�$�T�h���F#шG��������r�����$�T�I �F#шG�F���G������r�����$�T��F#шG�F�G�F���G�������V�������$�T�I  (08K�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�T��dl|��D$^_Ð�F�G�D$^_ÍI �F�G�F�G�D$^_Ð�F�G�F�G�F�G�D$^_Í�$    W�ƃ�����   �у���te��$    �fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tO������t��    fof�v�Ju��t*����t���v�Iu�ȃ�t��FGIu���    X^_Í�$    ���̺   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̋T$�L$��t�D$�%Ⱦs�L$W�|$��]�T$���   |�%��K�  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�Q�d蹝  Y�U��A	P�E��	P�A  ��Y�Y@]� U��V��������EtV���Y��^]� U���   �} t�d�  ��]ø��������v��������]��������������������������n��U��V�uW�����u��A  �    ��z  ��E�F�t9V��   V��藩  V�	�  P�'�  ����y�����~ t�v�  �f Y�f ��_^]�jh8q�&w  ����}�3��u������u�gA  �    �Rz  ���@w  ��F@t�f ��V�j  Y�e� V�?���Y���}��E������   �ǋu�}�V�  Y�U��V�u��u	V��   Y�/V�,   Y��t�����F @  tV�0�  P��  Y��Y��3�^]�U��SV�u3ۋF$<uB�F  t9W�>+~��~.W�vV��  YP脩  ��;�u�F��y����F��N ���_�N�f �^��[]�j�W   Y�jhXq��u  �u��u	V�<   Y�%V�h
  Y�e� V� ���Y���}��E������   ���v  Ëu�}�V�
  Y�jhxq�u  3��}�!}�j�@  Y!}�3��]�u�;5���   ������t]�@�tWPV�(
  YY�E�   �����@�t0��uP����Y���tG�}����u�@tP�n���Y���u	E܃e� �   F녋]�}�u���4�V�(
  YY��E������   ����t�E��$u  Ë]�}�j��  Y�jh�q��t  3��}�3��u������u�?  �    ��w  ����   V�	  Y�}��F@uqV�*�  Y�Ѓ��t���t���������������@$u)���t���t���������������B$�t�>  �    �mw  ����}��u�Nx
��8@��	V�P�  Y���}��E������   ���*t  Ëu�}�V��  Y�U��} u�">  �    �w  ���]�V�u��u�>  �    ��v  ���^]��u��  �#�Y�V���t�3���jh�q�us  3��}�3��u������u�=  �    �v  ����   V��  Y�}��F@uqV�ܣ  Y�Ѓ��t���t���������������@$u)���t���t���������������B$�t�4=  �    �v  ����}��u#�Nx��M�����V�u�;�  YY���}��E������   ����r  Ëu�}�V�s  Y�U��} u��<  �    �u  ���]ËE��t�j �p�0�u�   ��]�jh�q�;r  3��u������u�<  �    �mu  ����?�}��t
��t��u�V�  Y�e� W�u�uV�*   �����}��E������   ���r  Ëu�}�V�  Y�U��V�uW�F����   �}��t
��t��u{���S�F��uV�v�  �]؋E�Y3���E�]V�E������FY��y����F��t�t�   u�F   W�uSV��  YP��  ��#��[;�t3ɋ���{;  �    ���_^]�U��QQ�MSVW��t�]��t�u��u�L;  �    �7t  3�_^[�Ã} t���3���;�w؋����F  ��t�N��   �M�����   �V��  t6�F�E���t,��   ;�s�É]�P�u�6�;����E�)F��+�E�];�r^��tV�����Y����   �M��Å�t3����+E���]�P�uV�נ  YP�n�  �����tQ�M���;�w��U+�;�r=�M��(�EV� P茴  YY���t(�E�NK�M���3�A�M����-����E������N +���3��u�����jh r�o  �} t$�} t3��u������u��9  �    ��r  3���o  �V��  Y�e� V�u�u�u�Q��������}��E������
   ���ȋu�}�V�2  Y�U��Q3��E�9Et�E�P�u�[j  YY��u����ËE�VP�\�  �u����r  YY��^��jh r��n  3��}�3��u������u�59  �    � r  ����   �]��t	��t��@uׅ�t
��@t�M��M�A�=���w�����M�u�V�  Y�}�V����V譠  YY�f�����N��t���N�Fj[�8�E��u%�]S�J/  Y��u������}�� �N  ���   �N�]�^�F��~�E������   ���Mn  Ë}�u�V��  Y�U��EPj �u�uh���   ��]�U��� �e� V�uWj3�Y�}���u�8  �    ��p  ����;9Et�V�>  Y�����E�I   �u�u��M�;�w�E��u�E��u�uP�U��_^��U��SV�uW����F@uoV���  Y�Ȼ��;�t���t�у�����������B$u%;�t���t��������������A$�t�U7  �    �@p  ��_^[]Ë];�t��Fu�F�t��Fu��~ uV���  Y�;Fu	�~ u�@���F@�t	8t@�밈�F�F�����F���jh@r�~l  3��u������u��6  �    �o  ����)V��   Y�e� V�u�����YY���}��E������   ���rl  Ëu�}�V�  Yá�Vj^��u�   �;�}�ƣ�jP�,  YY����ujV�5��,  YY����ujX^�3ҹX���� �R��آ}����3�^������=�� t��  �5���   �%� YøX��U��V�u�X�;�r"����w��+�����P��  �N �  Y�
�F P�(�^]�U��E��}��P��  �EY�H �  ]ËE�� P�(�]�U��E�X�;�r=��w�`���+�����P��  Y]Ã� P�,�]�U��M�E��}�`����AP��  Y]Ã� P�,�]�U��j
j �u���  ��]�U��} t-�uj �5��P���uV��4  ���L�P��4  Y�^]������������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[�U��V�u��u3��m�E��u��3  j^�0��l  ���SW�}��t9urVWP�%�����3��6�uj P�c�������u	�3  j�9us�3  j"^�0�l  ���jX_^]�����SV�L$�T$�\$������tQ+���   t�
:uH��D�B��v4��u�
%�  =�  wً
;u҃�v����������#Ʃ����t�3�^[Íd$ ���^[�U��V�u���i   ����^]� U��V�EP���   ����^]� U��EV��f �p�F �0�   ��^]� U��E�p� �A�A ��]� U��V�u��f �p�F �   ��^]� �p�   U��VW�}��;�t�   � t�w���5   ��G�F_��^]� U��V���p�R   �EtV����Y��^]� U��} S��t-W�u�6  �xW�O  YY�C��t�uWP�e������C_[]� V��~ t	�v�����Y�f �F ^ËA��u�x�U��E�� VWjY���}��M_^��t� t��@��@�M��E���t� t�E� @��E�P�u��u��u��T��� U��V��u�N3�����j V�v�vj �u�v�u�6  �� ^]�U��QS��E�H3M�Q����E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u��  �� �E�x$ u�u�u�  j j j j j �E�Ph#  �|   ���E��]�c�k ��3�@[��U����H��e� �M�3��M�E��E�E�E@�E��.�M��E�d�    �E�E�d�    �uQ�u�\�  �ȋE�d�    ����XY�$��U���8S�}#  u��0�M�3�@�   �e� �E�/�H��M�3��EЋE�EԋE�E؋E�E܋E �E��e� �e� �e� �e�m�d�    �EȍE�d�    �E�   �E�E��E�E���v  ���   �E��E�P�E�0�U�YY�e� �}� td�    ��]ȉd�    �	�E�d�    �E�[��U��QQ�ES�]�HV�pW�M����u���x5�U���u��  �M��UN��k�9T};T~���u�}�K�u���y΋EF�0�E�8�E;xw;�v�L�  �M�k�_�1^[��U��QS�E���E�d�    �d�    �E�]�m��c���[�� U��QQSVWd�5    �u��E��1j �u�u��u�X��E�@����M�Ad�=    �]��;d�    _^[�� U��MV�u��u  ���   �N�u  ���   ��^]�U��V�~u  �u;��   u�nu  �N���   ^]��]u  ���   �	�A;�t�ȃy u�^]�I�  �F�A��U���/u  ���   ��t�M9t�@��u�3�@]�3�]�U���SVW��E�3�PPP�u��u�u�u�u�  �� �E�_^[�E���]�jh`r��b  �E��uz�V�  ��u3��F  ��u  ��u�R�  �����  �\����J�  ���&�  ��y�,v  ����  ��x ��  ��xj ��_  Y��u����   蛢  �Ʌ�ue����~�H���e� �=�� u�_  �|^  �u��u�c�  �u  趾  �E������   �   �u��u�=@��t�u  ��p��u^�5@���'  Y��u[h�  j�"  YY���������V�5@��'  YY��tj V�!t  YY�`���N��V����Y�������uj �<s  Y3�@��a  � U��}u�y�  �u�u�u�   ��]� jh�r�ea  3�@�u��u95���   �e� ��t��u5����t�uV�u�щE����   �uV�u�����E����   �]SV�u�/������}��u(��u$SP�u����SW�u���������tSW�u�Ѕ�t��u*SV�u�������#��}�t����tSV�u�Ћ��}��E��������&�M�Q�0�u�u�u�   ��Ëe��E�����3��`  �U��}u�uj �u�G����u�u�	�  YY]�U��V�u���woSW����u�\W  j�W  h�   �)\  ��YY��t���3�AQj P�d�����u&j[9,�tV�6�  Y��u���,*  ��%*  ���_[�V��  Y�*  �    3�^]������������̃=|� ��  ���\$�D$%�  =�  u�<$f�$f��f���d$���  � �~D$f(�f(�f(�fs�4f~�fT f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�q�  ���D$��~D$f��f(�f��=�  |!=2  �fT��\�f�L$�D$����f��fV�fT�f�\$�D$�U���uj �u�u�u�   ��]�U��� �e� Wj3�Y�}��9Eu�(  �    �a  ����x�EV�u��t��u�{(  �    �fa  ����S�����M�;�w�E��u�E��u�E�B   �u�u�P�u��8�  ������t�M�x�E��  ��E�Pj �T�  YY��^_��U���SVW�u3ۍM���]��������E��t9]t�9]t9]u��'  �    ��`  ��   �E�SSj��uS�p�D��E���u�L�P�'  �   �P�8  Y�E���tu�u�P�E�j��uS�p�D���tŋE�P�  ��Y��tI�u�u�u�u��uV�!2  ������t+�E�SS�u�uj�VS�p�@���u�L�P��&  ��YV�%����u�����YY�߀}� t�M��ap�_^��[��U��j j �u�u�u�u�������]�U��V��  ����t�uV�   ���Y��Y#�^]�U���SV3�W�}�]��]�]���u�&  j^�0�}_  ��_^[��j$h�   W�)����u����t�9^|9s�Y&  j^�0��jX9F|
�>�o@�w��g�  �E�P��  Y����  �E�P���  Y����  �E�P���  Y����  �^���|n���� vd�E��+ȍE�P�W�M�]����  YY���K���9E��<  W�=�  Y���-  �E��)E�E�PU�W��  YY�������G    �  VW��  YY�������9E�t-W���  Y��t"�E�E��G    ��ȋ���+�։U������؋E���+��j j<VS���  ���y��<��ĉ���j j<VS��  ���G�ڙj �j<�SV��  �G��y��<��ĉG���j j<SV���  ���G�ڙj �j�SV��  �G��y�����G���j jSV��  �ȅ�|+��t�G�j�^��O�WO3���������|��s�G����j^��O�G�W��у��G��m  G�O�G   �SSSSS�@]  �U��QQ�E�P�h��M��E�j �� ��*h��� !Nb�PQ��1  ��|=�o@�v����ЋM��t��Q�ú���  ��L�  ���������z�����������������̃��\$�D$%�  =�  ��   �<$�$������   f����%�  =�  t0��% �  u�Q����f�$�<$ uP�� �  uHf���� u>�ً���u$f��%��  uf��%��  uf�� %��  t�f�$�L$��  ��$    �D$  ���1   ���T$�ԃ��T$�T$�$��  fD$���f�$�O  �$�~$��Ë��L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�ËM�d�    Y__^[��]Q�Pd�5    �D$+d$SVW�(��H�3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(��H�3�P�e��u��E������E�d�    �U��V�u�<�� uV�q   Y��uj�sT  Y�4���(�^]�VW����S���t�tS�0�S�m����' Y���� �|�[�> t�~u�6�0����� �|�_^�jh�r��V  �=� u��M  j�FN  h�   �R  YY�}�<�� u[j�  Y����u��   �    3��Aj
����Y�e� �<�� uh�  V�l��4���V����Y�E������	   3�@�xV  �j
�7   Y�VW������~u�>h�  �6���l����� �|�3�_@^�U��E�4���,�]�jh0s��U  �E��tr�8csm�uj�xud�x �t�x!�t	�x"�uI�H��tB�Q��t'�e� R�p������E������%3�8E��Ëe�育  �t�@���t�Q�P�U  �U��V�u�������h��^]� �h� ���U��V���h�����EtV����Y��^]� j0h�r��T  �E�E�3ۉ]ȋ}�G��E؋u�v�E�P�����YY�E��f  ���   �E��f  ���   �E��f  ���   �{f  �M���   �]�3�@�E�E��u �u�u�uW�g������E�]��   �u���  YËe��4f  3ۉ��  �U�}�z�   �O��O�M��B�E�ÉE�9Bv?��k��z;L>�}~%�U;L�Uk��J�D@�E��J���M��	@�E�;Br�QRSW�	  ���]�]��u�E������E    �   ���T  Ë}�u�E؉G��u������Y�xe  �MЉ��   �je  �M̉��   �>csm�uH�~uB�~ �t�~!�t	�~"�u'�}�}� u!��t�v�����Y��t�uV�d���YY��}��j�.�������d  ���    t���  �e� �[�  ��d  �Mj j ���   �����U��}  W�}t�u �uW�u�  ���}, �uuW��u,����V�u$�6�u�uW�U  �Fh   �u(@�G�E�p�u�uW�u������,^��tWP�!���_]�U��E� �8csm�u9�xu3�x �t�x!�t	�x"�u�x u�d  3�A���  ��]�3�]�U���<�ESVW�}3ہ�   �]܈]��@��@�E����|;G|�Ԯ  �u�>csm���  �~�  �~ �t�~!�t�~"���   9^��   �c  9��   ��  �sc  ���   �hc  ���   jV�E�E���  YY��u�R�  �>csm�u+�~u%�~ �t�~!�t	�~"�u
9^u��  �c  9��   tl�c  ���   �E���b  �u쉘�   V�  YY��uD�}�9�  �É]�Oh ��L��������  �EC���E;|���  �E�E��E�>csm���  �~��  �~ �t�~!�t�~"��f  9_��   �E�P�E�P�u��u W�����M���;M���   �P�E��U�Z��]ԋ]9B���   ;B���   �:�}�z��}����}��   �M�F�@�P� �#�v�PQ�E��d  ����u*�E�U�M�H���E�U��ӋE�H���E��M����'�u��E��u$�u �u��u��u�W�u�uSV������,�U�E��M�A���M��U�;M��<���3ۀ} t
jV����YY�}� uy�%���=!�rk� te�wV��  YY��uV�+a  �&a  �!a  ���   �a  �}$ �M���   Vuz�u�x�E9_v8]u1�u$�u �u�W�uP�uV�s   �� ��`  9��   t�ҫ  _^[��� �  jV����YY�EP�M��Ep�^���h�s�E�P�E�h�v����u$����j�W�u�u�C  ���w�^����U��QQW�}�?  ��  SV�N`  ���    �]tHj �8����3`  9��   t1�?MOC�t)�?RCC�t!�u$�u S�u�u�uW�}���������   �{ u���  �E�P�E�P�u�u S�(����M��U���;�sy�p�E;F�|c;F�^��~���|��t�V�\�U��{ �]u8�~���ǋ}� @u(j�u$�N��u Qj PS�u�u�uW�����U��M���,�EA���M�;�r�^[_��U��QQSV�uW��tl3ۋ�9~]�ˉ]�E�@�@�P� �U��E���~5�E�p�F�2�P�  �M����u�E��U�H���E��U������G���M;>|�_^��[���ک  ��  ���^  3�9��   ���U��M�U�V�q�x�I��
��^]�jhs�L  �U�M�   �t����yz�e� �uVRQ�]S�W   ��HtHu4j�FP�s����YYP�vW������FP�s�s���YYP�vW�����E������L  �3�@Ëe��I�  �jh�s�(L  3ۋE�H���a  8Y�X  �H��u�    ��E  ��}��x����]�j��tB�u�v���  YY����   jW���  YY����   �N��E��PQ�����YY���   �u�E�p�tN��  YY����   jW��  YY����   �v�E�pW�������~��   �? ��   �FP�7�9^u9�V�  YY��tcjW�H�  YY��tU�v�FP�E�p�/���YYPW�M������:��  YY��t*jW��  YY��t�v��  Y��t�j [��C�]��誧  �E��������3�@Ëe��˧  3���J  �U��E� �8RCC�t!�8MOC�t�8csm�u*�\\  ���    钧  �K\  ���    ~�=\  ���   3�]�jh�r�UJ  �E�x�   �E�p��p�u��\  ���   �e� ;ut_���~�E;p|��  �M�A���U��E�   �|� t'�E�Ph  P�A�t��r�  ��u��)���YËe�e� �u��u���E������   ;ut荦  �E�p��I  Ëu��o[  ���    ~�a[  ���   �U��SVW�O[  �M�U3��csm�"�9��  u!9t�:&  �t�%���;�r
�A ��   �Bft!9q��   9uu}j�Q�u�u�������j9qu�%���=!�rW9qtR9u2�zr,9zv'�B�p��t�E$P�u �uQ�u�u�uR�փ� ��u �u�u$Q�u�u�uR������ 3�@_^[]�U��V�uW�F��tG�H�9 t?�}�W;�t�BPQ��  YY��t3��$�t�t�E� t�t�� t�t�3�@_^]��Z  �ЋBl;��t����Jpu��P  ���   �U����u�M������M��yt~�E�Pj�u�$�  ��������   �E�A���}� t�E��`p�����U����u�M������M��yt~�E�Pj�u���  ��������   �E�A���}� t�E��`p�����U����u�M��e����M��yt~�E�Pj�u��  ��������   �E�A���}� t�E��`p�����U����u�M������M��yt~�E�Pj�u�4�  ��������   �E�A���}� t�E��`p�����U����u�M�������M��yt~�E�Ph�   �u���  ��������   �E�A��   �}� t�E��`p�����U��=� u�M�P��H��]�j �u�C���YY]�U��=� u�M�P��H��]�j �u�h���YY]�U��=� u�M�P��H��]�j �u����YY]�U��=� u�M�P��H��]�j �u����YY]�U��=� u�M�P��H%�   ]�j �u�����YY]�U��} u3�]�SW�u�  �xjW�j�  �؃���t�uWS��  ����u
���3�_[]�3�PPPPP��H  ��.W  �ЋBl;��t����Jpu��M  �@��W  �ЋBl;��t����Jpu�M  �   �U���D�H�3ŉE�S3�V�u�]ԋ��   �]��]܉]�]؉u��]����  W�~9uWh  P�E�SP�>  ������  j�  jh�  �E��Q  jh�  �E��B  jh�  �E��3  jh  �E��$  �ȋEԃ�$�M؅��^  9]��U  ���M  9]��D  9]��;  ��È@=   |��E�P�7�p����  �E���  �M�S�7���EЋEܺ�   R�   PRAQh   ���   �M�S�I  ��$����  �E�S�7��   Q�   PQ�u�h   ���   S�  ��$����  �}�~18]�t,�}؍M���t�Q�����: �B;�~��8Y�uݍ~�E�S�7   Ph   �u�jS��  �����?  �}��E�3�f���   �M܃逈Y��X�考}���MĉEȈ~E8]�t@�M���t7�Q���;�$��   �P�E̋�� �  f��B�;�~�}���8Y�u�h�   ��   PW�{����M�j��   PQ�i����M�j��   PQ�W������   ��$��tHP�$���u=���   -�   P��������   ���P��������   ���P�������   �������E��    ���   ��   ���   ���   ���   �Eĉ��   �Eȉ��   �EЉFt�&�u��e����u��]����u��U����u��M���3ۃ�C�u��?���Y��_�D���   ��tP�$����   ���   ǆ�   �ǆ�   ǆ�   ��Ft   3��M�^3�[�*�����U��QQ�H�3ŉE�SV�uW��~!�E��I�8 t@��u������+�H;ƍp|���M$3���u�E� �@�E$��3�9E(j ��j V�u��   PQ�D��ȉM���u3��X  ~Kj�3�X���r?�M   ��   w���xT  �܅�t���  �Q������Y��t	���  ���M��3ۅ�t�QSV�uj�u$�D�����   �u�j j VS�u�u�6  ��������   �   �Mt,�M ����   ;���   Q�uVS�u�u��5  ���   ��~Bj�3�X����r6�}   ;�w�S  ���tf���  �P�������Y��tQ���  ���3���t@WV�u�S�u�u�q5  ����t!3�PP9E uPP��u �uWVP�u$�@���V蛿��YS蔿��Y�Ǎe�_^[�M�3��A�����U����u�M��t����u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap���U��VW3�j �u�u���  ������u'9H�vV�4����  ��;H�v������uË�_^]�U��SVW�=H�3��u������Y��u%��t!V�4��=H����  ��;�v������u�_^��[]�U��VW3��u�u�E�  ��YY��u,9Et'9H�vV�4����  ��;H�v������u���_^]�U��VW3��u�u�u��  ������u,9Et'9H�vV�4����  ��;H�v������u���_^]�j h t�>  3ۉ]���u��tph���VSS�E�P�Y�  ����t��t��"u
SSSSS�9A  j�u�����YY����u3��g  j�V�u�WS��  ����t��tă�"t���t	W����Y��W�uV�W  �؉]W���������t��FO  �E��Hl�MЋHh�M�3��}�E�PWSWW�E�P�7�  ����t��t��"u
WWWWW�V������e����E��P����Y���}܅��K����_�]؍E�Pj��u�u�Sj ���  ����t��t��"u3�PPPPP��������5����}�j�q���Y�e� ��D���tP�$���u
�t�����Y�E��@pu&���u�D���tP�$���u
�t������Y��M܉�L��\��E������   ���<  Ë]�j�U���Y�jh t�;<  �e� 3��}������u�~  �    �i?  3��~3��]������t�3�8����t���  ���u��u�C  �    �ȃe� �? u �-  �    j��E�PhH���  ���V�uSW�v�  �����}��E������   ����;  Ëu�}�V�v���Y�U��V�u�F��u��  �    ����nS�]���W�F��uV���  �}�Y3���}V������FY��y����F��t�t�   u�F   SWV�k  YP��  ��3Ƀ����_[�A�^]�jh@t��:  3��u������u�/  �    �>  ����<�}��t
��t��u�V�0���Y�e� W�uV���������}��E������   ����:  Ëu�}�V�h���Y�U�졠�3H�t�u��]�]�%��U�졤�3H��ut��]����]�U�졨�3H��ut��]����]�U�졬�3H��u�ut��]����]�U�조�3H�t�u�u�u��]��u�u�l�3�@]�U��QV�5(���y%��3�3H��u�tV�M�Q�Ѓ�zuF�5(�3�����^��VWh�����5����h�W��3H�h�W�����3H�h�W�����3H�h�W�����3H�h�W�����3H�h�W�����3H�h W�����3H�hW�����3H�h0W�����3H�hDW�����3H�hdW�����3H�h|W�����3H�h�W�����3H�h�W�����3H�h�W�����3H����h�W��3H�h�W�����3H�hW�����3H�h4W�����3H�hHW�����3H�hdW�����3H�hxW�����3H�h�W�����3H�h�W�����3H�h�W�����3H�h�W� ���3H�h�W����3H�h�W����3H�h�W����3H�_��^�U���u���P���]�U��j �x��u�t�]�U��U�,��M#M��#�щ,�]��L�  ��tj�j�  Y�,�t!j�a ��tjY�)jh  @j�8  ��j�4  ���������������̋T$�L$��   u@�:u2��t&:au)��t��:Au��t:au������uҋ�3���������Ë���   t���:u����t���   t�f���:u΄�t�:auń�t��������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^���G  ��u���Ã��U��V������MQ��    Y���   �0^]��G  ��u���Ã��U��M3�;Ő�t'@��-r�A��wjX]Í�D���jY;��#���]ËŔ�]�U���V�u�M��3����u�E�M�L0u3�9Ut�E����   �p#E���t3�B�}� ^t�M��ap�����U��jj �uj ������]�U��Ef���f��u�+E��H]�U���ESVW��Y�9  ��  ��I��   ��   ����  ��	��  ����   ��t`Ht1���  �E�@���a  ���X  �u �u�ujP�V  �E�H���9  ���0  �u�E�u���  �J  �E�H���  ���  �u�E�u����   �  �Mj%�Zf��E���  �E�@����  ����  j�Y����u���u �u�ujR�  ��M��   jY+���   HHtPHHt-H��  �u�u�u�uj�u�  ������  �j  �U�B���L  ;��D  ��t�H���U�B���-  ;��%  �ȋB���  =m  �  ;�}3�����j�^��;������@�����E�8 ��  �8;��  �u �u�uj�0��   �E�@����  ��;�S����E�@=������  =�  ��  jd�Y���u �u�uj��k�d��*�����m��  �U  ��Z��  ���  H��   HthHt3���P  �E�@���2  =m  �'  �u @�u�uj������E�x�	  �x��   �u �u�uj�p�6  ���  �}  �ut@�u�}VW�uj�u�  ������   �> ��   �j Y�uf���VW�$����}�]WS�u3�V�u��  ������   97��   �j Y�uf���WS������E�H��xQ��L�u�E�u����   �f  �E�H��x-��(�u�E�u����   �B  �E�@��x	�������_����    �J4  3�_^[]Ã�p��   ����   H��   Ht[Hu��U�  �u3�j��u虤  �M�}�]3�9q ���4��E�7�3P�(�  ������   �M�M����3�@+��   �E�@���d����u ��u�ujjdY�������}  �u�u�u�utj�����j �����E�@��� ����������u �u�uj�����E�@���������������u�u���E��L  �	�M��P  ��   ��3�@�����VVVVV�!3  �U��V3�9ut�u�u�u�V   ���N�M�E;sBHS�XW�}��t*� �E��E
   �}�E���0f��EF�I�KuߋM�6)1_[��1^]�U��MV�1W�}�?v#S�]�Ùj
[���؍B0f������~�?w�[��1���f�f�f�
����;�r�_^]�U��M�9 t!�UV�uW�:f��t���f�8��	u�_^]�U���0�H�3ŉE��E�U�M�EЋE�E��ES�]V�E؋�3�W�UԉM�+�tHt��\  ���X  ���T  ���   �)  ����۸l  fBVf�E�f�Bf@f�E�f�Bf�E�f�Bf�E�f�Bf�E�f�f�E�3�VWf�E��E�P��V��`  ��t�#  ��"  ���E����   �E   =   w�A  ��u����   ���  �P������Y�u��t���  ���u��to�u�E�VWP�E�j ��`  ��t�"  ��"  �Ѓ�J����~#�]؋u��; v�f�f�����J���u�V�E���Y3�@�e�_^[�M�3��������7f��t�]؃; tۃe� 3ɋ��փ�A�;�t��]�]؃�d�  ��   j'X;���   ��At��HtP��Mt��a��  hW��  YY��uJ��
�^ItItItI��  jB�  jb�  �E�   jm�  ItIt�q  �E�   jH�~  hW�I�  YY��u����}�jp�a  �<O���s  �f��������U��; �[  ��f;��O  �j'f����Xf��u��5  ItItItI��   jA��   ja��   �E�   jd��   ��h��   ����   ����   Jt#����   IItII��   jY�   jy�   �Eԃx�E���L  ���P  ��u�; v�u�f��f����%�
f��t�u��; v���f����
f��u�}��hItIt	�$�E�   jS�4ItIt	��E�   jM�!ItIt�U����f�0���*�E�   jI�}�X�u��u�S�u��u�P�u��$�������t�7f�����������3��~���U����ESVW�u�M�3��E�詨���E����   �]����   �}3�f�����   �U��u�E䋐�   �U�ÉE�����   �M��]��ۅۋ]tn�]�f��%�]t�E�f��M�E�����H�M�E��@9ut|����f�?#u3�@��PR�E�P�EP��uP�E�P�9�������t �M�E����U��u���t3���f�+u��:9u�v3�@��ƋM�3�f���u9U�w����� "   ��
����    ��,  �}� t�M�ap�_��^[��U����M�SW�u�q����]�   ;�s`�M�yt~�E�PjS膭  �M������   �X����t�}� ���   �t�E��`p�����   �}� t�M��ap����   �E�xt~-�����E�M���QP�+�  YY��t�Ej�E��]��E� Y��1���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QW���   �E�P������$��u8E��{����E��`p��o�����u�}� �E�t%�M��ap���U��E���Ѐ}� t�M��ap���_[��U��=� u�M�A���w�� ��]�j �u����YY]����̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� U��S�]��V�� ��  H��  H��  H�=  �UH��  �uW�� ��  �;��   ���+�t3Ʌ����M��������  �~�B+�t3Ʌ����M�������y  �~�B+�t3Ʌ����M�������W  �N�B+�t3������E�����3Ʌ��1  �F;Bt���B+�t�����M�������
  �~�B+�t3Ʌ����M��������  �~�B+�t3Ʌ����M��������  �N�B+�t3������E�����3Ʌ���  �F;Bt���B+�t�����M�������y  �~	�B	+�t3Ʌ����M�������W  �~
�B
+�t3Ʌ����M�������5  �N�B+�t3������E�����3Ʌ��  �F;Bt���B+�t�����M��������  �~�B+�t3Ʌ����M��������  �~�B+�t3Ʌ����M��������  �N�B+�t3������E�����3Ʌ��~  �F;B��   �B�~+�t�����M�������R  �~�B+�t3Ʌ����M�������0  �~�B+�t3Ʌ����M�������  �N�B+�t3������E�����3Ʌ���  �F;Bt���B+�t�����M��������  �~�B+�t3Ʌ����M��������  �~�B+�t3Ʌ����M�������}  �N�B+�t3������E�����3Ʌ��W  �F;Bt���B+�t�����M�������0  �~�B+�t3Ʌ����M�������  �~�B+�t3Ʌ����M��������  �N�B+�t3������E�����3Ʌ���  �F;Bt���B+�t�����M��������  �~�B+�t3Ʌ����M�������}  �~�B+�t3Ʌ����M�������[  �N�B+�t3������E�����3Ʌ��5  j Y+���;��_����Ӄ��  �$�@��F�;B���   ���B�+�t3Ʌ����M��������  �~��B�+�t3Ʌ����M��������  �~��B�+�t3Ʌ����M��������  �N��B�+�t3������E�����3Ʌ��y  �F�;B���   ���B�+�t3Ʌ����M�������L  �~��B�+�t3Ʌ����M�������*  �~��B�+�t3Ʌ����M�������  �N��B�+�t3������E�����3Ʌ���  �F�;B���   ���B�+�t3Ʌ����M��������  �~��B�+�t3Ʌ����M��������  �~��B�+�t3Ʌ����M�������q  �N��B�+�t3������E�����3Ʌ��K  �F�;B���   ���B�+�t3Ʌ����M�������  �~��B�+�t3Ʌ����M��������  �~��B�+�t3Ʌ����M��������  �N��B�+�t3������E�����3Ʌ���  �F�;B���   �B��~�+�t3Ʌ����M��������  �~��B�+�t3Ʌ����M�������d  �~��B�+�t3Ʌ����M�������B  �N��B�+�t3������E�����3Ʌ��  �F�;B���   ���B�+�t3Ʌ����M��������   �~��B�+�t3Ʌ����M��������   �~��B�+�t3Ʌ����M��������   �N��B�+�t3������E�����3Ʌ���   �F�;B�tu���B�+�t3Ʌ����M������u`�~��B�+�t3Ʌ����M������uB�~��B�+�t3Ʌ����M������u$�N��B�+�t3������E�����3Ʌ�u3ɋ�_��  �F�;B�tu���B�+�t3Ʌ����M������u��~��B�+�t3Ʌ����M������u��~��B�+�t3Ʌ����M������u��N��B�+�t3������E�����3Ʌ��q����F�;B���   ���B�+�t3Ʌ����M�������D����~��B�+�t3Ʌ����M�������"����~��B�+�t3Ʌ����M������� ����N��B�+�t3������E�����3Ʌ�������F�;B���   ���B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M�������i����N��B�+�t3������E�����3Ʌ��C����F�;B���   ���B�+�t3Ʌ����M�����������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ�������F�;B���   ���B�+�t3Ʌ����M�����������~��B�+�t3Ʌ����M�������]����~��B�+�t3Ʌ����M�������;����N��B�+�t3������E�����3Ʌ������F�;B���   �B��~�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ��}����F�;B���   ���B�+�t3Ʌ����M�������P����~��B�+�t3Ʌ����M�������.����~��B�+�t3Ʌ����M�����������N��B�+�t3������E�����3Ʌ�������B��N�+������3������E����������F�;B���   ���B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M�������t����~��B�+�t3Ʌ����M�������R����N��B�+�t3������E�����3Ʌ��,����F�;B���   ���B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ�������F�;B���   ���B�+�t3Ʌ����M�������h����~��B�+�t3Ʌ����M�������F����~��B�+�t3Ʌ����M�������$����N��B�+�t3������E�����3Ʌ�������F�;B���   ���B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ��g����F�;B���   ���B�+�t3Ʌ����M�������:����~��B�+�t3Ʌ����M�����������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ�������F�;B���   �B��~�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M�������^����N��B�+�t3������E�����3Ʌ��8����F�;B���   ���B�+�t3Ʌ����M�����������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ������f�F�f;B�������D  �F�;B���   ���B�+�t3Ʌ����M�������a����~��B�+�t3Ʌ����M�������?����~��B�+�t3Ʌ����M�����������N��B�+�t3������E�����3Ʌ�������F�;B���   ���B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ��`����F�;B���   ���B�+�t3Ʌ����M�������3����~��B�+�t3Ʌ����M�����������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ�������F�;B���   ���B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M�������z����~��B�+�t3Ʌ����M�������X����N��B�+�t3������E�����3Ʌ��2����F�;B���   �B��~�+�t3Ʌ����M�����������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ�������F�;B���   ���B�+�t3Ʌ����M�������m����~��B�+�t3Ʌ����M�������K����~��B�+�t3Ʌ����M�������)����N��B�+�t3������E�����3Ʌ������F�;B���   ���B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������~��B�+�t3Ʌ����M������������N��B�+�t3������E�����3Ʌ��l����~��B�+�t3Ʌ����M�������J����B��~�+��T���3Ʌ����M�����9����M��1+�t3������E��������   �q�B+�t3������E��������   �q�B+�t3������E��������   �I�B+�t3������E�������   �U�u�
�+�t3������E������uj�J�F+�t3������E������uL�J�F띋U�u�
�+�t3������E������u �J�F�n����E��E� �]���3�^[]ÍI Jwf{����v�zI�0v7z|~���u�y�}�u	yN}��jtrx�|��s�w |U�<sTw�{�U���,�H�3ŉE��E�MS�E��EV�u�EԋEW�E�M܅�~"VP�2  YY�M܋��} ��~WQ�  YY������}�3���  ���|�E$3ۉ]؅�u�E�� �@�E$��t����   ;�ujX��  ��~3�@�  ��~j��M�QP�p���t���~+�}�r�E�8]�tۋu�H��tъ:r:�v���8u�뾅�~2�}�r��E�8]�t��u܊H��t��:r:��z�����8u��{���SSV�u�j	�u$�D��ȉM�������~Ij�3�X���r=�M   ��   w���@"  �܅�t���  �Q�N�����Y��t	���  ���M��������QSV�u�u$jV�D�����   3�PPW�u�j	V�D��ȉM����   ~Kj�3�X���r?�M   ��   w���!  ���t���  �Q�í����Y��t	���  ���M��3���t5QVW�u�j�u$�D���t�u�V�u�S�u�u��  ���E�V蟍��YS蘍���E�Y�e�_^[�M�3��D�����U��E�U�ȅ�tI�: tB��u�I+�H]�U����u�M��W����u$�E��u �u�u�u�u�uP�F����� �}� t�M��ap���U��V3ɾ�   ��+U��+� t��y�p���H;�~܃��^]�U��SVW3���   �;�+���jU�4�@�u�  ����ty�^���~;�~Ѓ�����D_^[]�U����3H�t3�QQQ�u�u�u�u�u�u��]��u�u�u�u�u�u�   YP���]�U��ESVW��t[=   tT=   tM�} �uu��@��x<P�����Y��x1��$jUS蝰  YY����~;�}SV�u��  ����u�G�3�_^[]�3�PPPPP�J  �U��} t�u�����Y��x=�   s	�� ]�3�]�U��j j �u�T�]� U����3H�tj �u�u�u��]ËEjh��T�����%T� ]�U����3H�tj �u�u�u�u�u�u��]��u�u�u�u�u�u�F���YP���]�U���u���3H��u�u�ut��]�����YP���]�U���u� �3H��u�u�u�u�ut��]������YP���]�U���3H��u�ut��]����P�6�����]�U���3H�t�u��]�j�u����YP���]�U���3H�t3�QQQ�u�u�u�u�u�u��]��u�u�u�u�u�u�@���YP���]�U��V�u3���t^�MSW�}jA[jZZ+��U�jZZ�f;�rf;�w�� ������f;�rf;Ew�� ����Nt
f��tf;�t�����_+�[^]�U��E��~P�u��  YY�u�uP�u�u�u������]��̃��$���  �   ��ÍT$訮  R��<$�D$tQf�<$t�`�  �   �u���=� �Ӯ  �   � ��Ю  �  �u,��� u%�|$ u���5�  �"��� u�|$ u�%   �t����-�C�   �=� �v�  �   � ���  Z�j�u�  Y��tj�h�  Y��u�=X�uh�   �1   h�   �'   YY�U��M3�;�X:t
@��r�3�]Ë�\:]�U����  �H�3ŉE�V�uWV������Y���y  Sj��  Y���  j�ݯ  Y��u�=X���   ���   �A  hl;h  h`���  ��3ۅ��/  h  h��Sf��������  ��uh�;Vh���Ό  ������   h������@Y��<v5h�������E���-��j��h�;+�VQ�j�  ������   h�;h  �`�V�ޭ  ������   Wh  V�ǭ  ����u{h  h�;V��  ���Wj��������tI���tD3ۋˊO�����f9Ot	A���  r�S�����P�����P�]��x���YP�����PV���[�M�_3�^�h�����SSSSS�
  �U���   �H�3ŉE��E�U�MSVW�}��l�����t������  h�   ��|�����P�u3�QR��p���諱  ����x�����ut�L���z��   VV�u��t�����l����y�  ����x�����tcjP�������YY��tS��x���ǅp���   S�u��t�����l����7�  ����x�����tjP������YY���u!9�p���tS�"���Y����M�_^3�[�R����Ë�x����A�PSQR�i�  ������   9�p���tS����Y3�����uN3�VV�u�7Q�:����؃���t'jS� ���YY���tSP�u��t�����������u��7蔚��Y�7�k������c���!�x���j��x���P�E    PQ����������:�����x�����k���VVVVV�8  �U��E���]�U��QS3�V9]u����j^�0��  ���   �u��t��������u�����u3�C3�PPj��u�PS�D��E���u�L�P����Y3��A�P�S���Y���t��u�Pj��uj S�D���u�L�P�g����6蓙���& Y�3�@^[��U��Q�E�Ph,<j �����thD<�u������t�u����U���u�����Y�u����VW�5���<��5������t�> t�6����Y��u�5��SV�����5��3�Y�����t9t�6����Y��u�5��V�՘���5������Ę���5��蹘�������������t9��tW藘��Yj��8�����$���tP�z���Y�$��(���tP�d���Y�(��5 ��$�[��u� �� �;�tP�8���Y�5 �_^�U��������u�I���Yh�   �   �jj j �1  ���U��=h thh�a�  Y��t
�u�hY��2  h��h����   YY��uPVWh���"w��Y�X��������t�Ѓ�;�r�=�� _^th�����  Y��tj jj ���3�]�U��j j�u�   ��]�Vj �8���V�_e  V��  V�����V蠮  V�%�  V�_  ��^�/���U��V�u����t�Ѓ�;ur�^]�U��V�u3����u���t�у�;ur�^]�j����Y�j�x���Y�jh`t�^  j�����Y�e� �=����   ���   �E����} ��   �5���5<��֋؉]ԅ�tt�5���֋��]�}��}܃��}�;�rWj �8�9t�;�rG�7�֋�j �8�����5���5<��։E��5���֋M�9M�u9E�t��M�ى]ԉE����h��h�������YYh��h�������YY�E������    �} u)���   j�e���Y�u�h����} tj�O���Y��   �U��} u�����    �r  ���]��uj �5����]�����������h �d�5    �D$�l$�l$+�SVW�H�1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q��������U���S�]VW�{3=H��E� �E�   ��s���t�O�30�����O�G�30�����E�@f��   �E�E�E�E�C��C�E������   �@�@�L������E���t{���R�  ��M����~   ~h�E�8csm�u(�=` th`�ê  ����tj�u�`���U�M�5�  �E�U�9PthH�V���6�  �E�X����tu�f�M��É]�����]�����tG�!�E�    ��{�t6hH�V�˺������  ����t�O�30��~���O�W�32��~���E�_^[��]ËO�30��~���O�G�30��~���M��֋I�e�  �U���(  �H�3ŉE��}�Wt	�u�Ǫ  Y������ jL������j P������������������0�����������������������������������������������f������f������f������f������f������f��������������E�������E������ǅ0���  �@��������E�������E�������E����������������P�����Y��u��u�}�t	�u�ԩ  Y�M�3�_�}����U��E���]�U���5���<���t]���u�u�u�u�u�   �3�PPPPP��������j�& ��tjY�)Vj� �Vj�u���V�.�����^�U��%ľ ��S3�C	�j
�}& ���  3ɋÉľ�V�5�W�}�����_�O�W�E�   �5�t���ľ   �5��E�   t���ľ   �5�j3�X��u���^�N�V�E�   �5Ⱦt	���5Ⱦ3�3���}���_�O�W�}�Genuu_�}�ineIuV�}�nteluM3�@3����_�O�W�E�%�?�=� t#=` t=p t=P t=` t=p u	���5Ⱦ_^3�[�������������̃=ľr_�D$�����fn��p� ۋT$�   ���#���+��o
f��ft�ft�f��f��#�u����������f~�3�:E��3��D$S�����T$��   t�
��:�tY��tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u!% �t�% u��   �u�^_[3�ÍB�[ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[�U��3�9Ev�M�9 t@A;Er�]�U��SV�5 �W�}W�փx t�wx�֋��   ��tP�փ| t�w|�֋��   ��tP��jX�_�E�{�P�t�; t�3�֋E�{� t�{� t�s��֋E��H�Eu΋��   �   P��_^[]�U��SV�u3ۋ��   W��tf=8�t_�Fx��tX9uT���   ��t9uP苎�����   ���  YY�F|��t9uP�m������   �z�  YY�vx�X������   �M���YY���   ��tD9u@���   -�   P�,������   ��   +�P�������   +�P�������   � ��������   =X�t9��   uP�i�  ���   �׍��YYjX���   �~�E��P�t���t�8 uP謍���3襍��YY�E�� t�G���t�8 uP舍��Y�E����H�Eu�V�r���Y_^[]�U��V�u����   SW�=$�V�׃~x t�vx�׋��   ��tP�׃~| t�v|�׋��   ��tP��jX�^�E�{�P�t�; t�3�׋E�{� t�{� t�s��׋E��H�Eu΋��   ���   Q��_[��^]�jh�t�Y����&	  ������Npt"�~l t�	  �pl��uj �l���Y���k����j�Ɵ��Y�e� �5���FlP�!   YY���u��E������   뼋u�j�����Y�U��W�}��t;�E��t4V�0;�t(W�8�����Y��tV�����> Yu����tV�O���Y��^�3�_]Ã=�� uj��P  Y���   3��U��E-�  t&��t��tHt3�]á`<]á\<]áX<]áT<]�U����M�j �)t���E�%� ���u��   ����,���u��   �������u�E���   �@�}� t�M��ap���U��S�]VWh  3��sWV��|��3��ȉ{�{��  ������{���� ���+��  �7�FIu���  �   �9�AJu�_^[]�U���   �H�3ŉE�SV�uW������P�v�p�3ۿ   ����   �È�����@;�r�����ƅ���� ��������Q���;�sƄ���� @;�v�����u�S�v������PW������PjS�6{  S�v������WPW������PW��  S�%�����@������S�vWPW������Ph   ��  S�������$����M�����t�L��������t�L ��������  ���  A;�r��Wj���  X+ˉ������������� ��w
�L�A �������w�L �A����������A��  ;�r��M�_^3�[�t����jh�t������  ������Opt�l t�wh��uj �����Y��������j�I���Y�e� �wh�u�;5 �t6��tV�$���u�� �tV�݈��Y� ��Gh�5 ��u�V� ��E������   뎋u�j�L���Y�jh�t�2��������  �؉]��=����sh�u�����Y�E;F�n  h   �����Y�؅��[  ��   �E�ph���3��3S�u�G  YY���}���  �E��ph�$����E�u�Hh�� �t
Q����Y�E�XhS� ��E��@p��   �����   j����Y�u��C�о�C�Ծ��  �̾�ΉM���}f�DKf�MؾA��ΉM���  }�D���A��u���   }��  �� �F���5 ��$���u� �= �tP�Q���Y� �S� ��E������   �1�}j�˛��Y��#���u�� �tS����Y������    �3���������U��� �H�3ŉE�SV�u�u�-�����Y�]���uV����Y3��  W3��ωM��9�(���   A��0�M�=�   r����  ��   ����  ��   ��P�������   �E�PS�p�����   h  �FWP��w���^3�C����  9]�vO�}� �E�t!�P��t�����LA;�v����8 uߍF��   �@Iu��v��������  �^��~3��ȋ�����~����   9=�tV�����   ����   h  �FWP�Tw���U��k�0��8��E�8 ��t5�A��t+������   s��$�D�AC;�v���9 u΋E�G���E��r��]�S�^�F   �W�������  j�N��,�_f�f��R�IOu�V�<���Y3�_�M�^3�[�Jp����jh�t�����u���   �~$ t	�v$����Y�~, t	�v,�ӄ��Y�~4 t	�v4�Ą��Y�~< t	�v<资��Y�~@ t	�v@覄��Y�~D t	�vD藄��Y�~H t	�vH舄��Y�~\8At	�v\�v���Yj誗��Y�e� �~h��tW�$���u�� �tW�I���Y�E������W   j�q���Y�E�   �~l��t#W����Y;=��t����t�? uW�>���Y�E������   V����Y������ �uj�~���YËuj�r���Y�U��@����t'V�u��uP������@�Yj P� ���YYV����^]�V�   ����uj�Y���Y��^�VW�L��5@����ɳ����Y��uGh�  j蠮����YY��t3V�5@������YY��tj V�%   YY�`��N���	V�"���Y3�W�|�_��^�jhu�����u�F\8A�f 3�G�~�~pjCXf���   f���  �Fh ����   j����Y�e� �vh� ��E������>   j����Y�}��E�Fl��u����Fl�vl�5���Y�E������   �R����3�G�uj����Y�j����Y�������������u�c   3��h%��_���Y�@����t�Vh�  j�n�����YY��t-V�5@�菲��YY��tj V�����YY�`��N��3�@^��   3�^á@����tP�����@��Y�=����Q�L$+ȃ����Y�*�  Q�L$+ȃ����Y��  jhhu�(������95��t*j輔��Y�e� Vh������YY����E������   �1����j����Y�3��U��} u3�]�SjU�u�E�  ��YY��Ur3���]   WP訬����Y��u_[]ÍCP�uPW苒  ����u����3�PPPPP������U��VW�}W�u�u�}p  ��3���uF���   f90tPhAj�u�u�~  ����   f97tWh Aj�u�u�]  ��_^]�VVVVV�n����U��QSVW�}h�  3�SW�r���u���f��u3���   j.Yf;�u-�Ff9t%jP��   jP跑  ������   f��  �ĉ]hAV��  YY����   �F�M���Mj,Z��u��@��   j.Yf;�tyPVj@W�:��u��@sh��_tcPVj@���   ���uR��sMf��tf;�uCPVj��   P�!�  ����u#j,Xf;��/���f���&����u����E�W���3�PPPPP����_^[��SSSSS�D����U��V�u��t�E��t;�tWj.Y���  P�����Y_^]�U����  �H�3ŉE��ES�]V�uW�}�����������V������   ��(������   �� ������  ��,���3ɉ�$�����u3��M�_^3�[��i�����  jUP�u�����S�$�  �����R  f�>Cu/f9Fu)�����hA�uV�n  �����'  ��t����V� ���Y�����=�   s,V��,����ר  YY����  V�� ������  YY����  �=��3=H���0������V��P���}���YY��uw��0���P����(���WPt�ݶ  ����  ����tW��0���P��   W��,��������������   ��P���P�I���@P��P���P�uS��  ������   �>  ��(���V�k���Y���  j��$���Ph  V��������t
��$�����u�����$�����������GWVh�   ��,���衎  ������   WV�uS苎  ������   WVjU������q�  ������   ��   3�f9t'�����;�s@PVW�� ����A�  ����tSSSSS�s�� ���3�f��������tj��(���W��g������,��������S�uV�l  ����u)������S����@PSjU������Ӎ  ����u�{���3�PPPPP�#����U��S3�V��9]~"W�}��7�u�u�,�  ����uF;u|�_^[]�SSSSS������jh0u�w���3ۉ]�}v������    ����3��>  �"������u�������Np!]�jh�   ����YY���}܅���   j�Ŏ��Y�E�   �vlW�)���YY�e� �   �u�uW�c  ���؉]����   �} thP��u�ݥ  YY��t
��   j�c���Y�E�   �FlWP�����W�������Fpu<���u3�vlh������YY������   �0����   � ��At����e� �   �.�}܋u�j�R���YË]�u�j�C���Y��W�-���W�����YY�E������   ���W���Ë]�u��fp��U���SW3�Gh�  �}�������3�Y����   V�sf��;�}�w$hA�5�?jhQ  V�������?�E��G$���E�hAhQ  V�%�  ������   �E�p�6�0芤  �����!E��E��΃��1�shA�0�M�jhQ  V�E������E��� =�?|��}� uM� t�w�$���u	�w�y��Y� t�w�$���u	�w�qy��Y3ɉO�O�_�w��^_[��S�Uy��� �5$�Yt�w�օ�u	�w�7y��Y� t�w�օ�u	�w�y��Y�G43ɉO�O�O�O�3�QQQQQ������U����  �H�3ŉE��ESV�uW�}��4�����t��tVPW�R  ���)  ��D��  3���ǅ@���   ��<�������  f�>L�^  f�~C�S  f�~_�H  h AV�ѣ  YY��8������&  ��+�����D����  j;Yf9�  ��D���ǅ@���   ��?WV�3�O�  ����u�3�í��Y;�t��@��������?~Ӌ�8�����hAV�Ȣ  ��4�����<���YY��D�����uj;Yf9��   ��@���bPV������h�   P�7�  �����  ��D����=  �  3�f������������P��@���W��   ������D���tC��<����4F3�f9t��f9���������   �   3��   PjU��H���Ph�   ������PV���������tw�G3���D�����t@�0������P葡  YY��t%������PVW�g   ������D���u3ɉ�@������D���C��@���F����D�����~���u���f���W�'���Y�M�_^3�[��a������  3�PPPPP�l����U����  �H�3ŉE�S�]V�uW�}��4��������  ��@�����,���PjU��H���Ph�   ������PV���������u3��M�_^3�[�Ka�������������t;�����P莠  YY��u�D;�̍�����P腫���p�u   Q�W���YY��$�����t��H�D;�� �����4�����(��0�������<���� ������G�����������PVQ�!e  ��3�����  f������C��0����D;uf9�����u
��<����1���H���P�����Y��<������4������u  ��,����G��@�����8����H ��(����H$��0����Ή�D�����8����G;��4�����   ��8�����8������(����I��8������0�����0�����D���A�Z�������4�����(�����D�����|���D�����@�������   j�w������Pjh�@jV�He  ������   �ƹ�  f!�E����@��r�h�   �5��������P�;�����@��������@�A�O��t���@�����D�����(��������D����D��A��D�������0����\�������L�����@����q�G��4�����A�Gp���u��,����G���u	��,����Gk�W���?���� ���Yt5�D;��<����3�fs����������$���P�Rs�������YY�G�)���=P�t<�t;�$���u.�t;�$s���t;�s����<����0�s����<����t;���0��$����    �D;����VVVVV������U����j���<�  �u�����=� YYuj�"�  Yh	 �����Y]�U���$  j�L ��tjY�)���������5��=ܿf��f���f�ؿf�Կf�%пf�-̿�� ��E ����E����E���������@�  ��������	 ����   � �   jXk� ǀ�   jXk� �H��L�jX�� �L��L�h$A�������U��j�   ]�U���  j�G ��t�M�)���������5��=ܿf��f���f�ؿf�Կf�%пf�-̿�� ��E ����E����E����������������	 ����   � �   jXk� �M���h$A������Å�uf���fn�f`�fa�fp� SQ�ك���ux�ڃ���t0ffAfA fA0fA@fAPfA`fAp���   KuЅ�t7����t��I f�IKu���t����t
f~�IJu���t�AKu�X[��ۃ�+�R�Ӄ�t�AJu���t
f~�IKu�Z�^���jh�u����j�0���Y�e� �u�F��t0�����M��t9u,�A�BQ��o��Y�v�o��Y�f �E������
   �}���Ë���j�8���Y�U��j �u�u�u�u�u�u�   ��]�U��E��et_��EtZ��fu�u �u�u�u�u��  ��]Ã�at��At�u �u�u�u�u�u�s  �0�u �u�u�u�u�u�   ��u �u�u�u�u�u��  ��]�U���,SVWj0X�u�ȉM��M��E��  3��QW���}��y���u��t�M��u	蜣��j��G�;�w芣��j"_�8�v�����  �U��Z�E����%�  =�  uy3�;�uu���;�t�A�j WP�^SR�  ������t� �  �;-u�-F�}j0X�������$�x�F�FjeP�<�  YY��t�����ɀ����p��@ 3��O  3���   ��t�-F�} �]j0X�����$�x��ۈF�J�����'��  �3���]�u'j0X�F�B�
%�� ���u3��E���E��  ��F1����F�M��u� ��Eԋ��   � � ��B%�� �E�w	�: ��   �e �E��   �M��~S��R#E#ыM��Ɂ��� 舭  j0Yf�����9vËM�U��E���E�E�����FO�M�E�f��y�f��xW��R#E#ыM��Ɂ��� �0�  f��v6j0�F�[���ft��Fu�H��]�;E�t���9u��:��	�����@���~Wj0XPV�%^������E�8 u���} �U����$�p���R�4踬  ��3��ځ��  #�+M��x;�r	�F+����F-������ۋ��0;�|A��  ;�rPRSQ芫  0�F3��U�;�u;�|��drPjdSQ�g�  0�F�U�3�;�u;�|��
rPj
SQ�D�  0��U�F�]�3���0��F���}� t�M܃ap���_^[��U��j �u�u�u�u�u�T  ��]�U����M�SW�u ��S���]��t�} w	�@���j��U3����ǃ�	9Ew�"���j"_�8������   �} t �M3�����P3��9-���P��  �UYY�EV�8-��u�-�s��~�F��E�F���   � � �3�8E�������9Et��+�Eh,APV�-J������ut�N9}t�E�U�B�80t-�RJy���F-jd[;�|��� Fj
[;�|��� F V�h�^t�90uj�APQ�J�����}� t�M��ap���_[��WWWWW�����U���,�H�3ŉE��ES�]VW�}j^V�M�Q�M�Q�p�0�ߨ  ����u�؞���0��������t�u��u
�����j^����;�t3��}�-����+�3�����+ȍE�P�CPQ3Ƀ}�-��3�������P��  ����t� ��u�E�j P�uSVW��������M�_^3�[�T����U����ES�@V�uH�M�E���Q���u��t�} w����j[������   3�W�}8]t�M�;�u�U3��:-���f�00 �E�8-u�-F�@��jV�  Y�0YF����~JjV�  �E�Y���   Y� � ��EF�@��y&8]t�������;�|��WV�`  Wj0V�-Z����_�}� t�M�ap�^��[��U���,�H�3ŉE��ESW�}j[S�M�Q�M�Q�p�0�-�  ����u�&�����������lV�u��u�������������S���;�t3��}�-����+ȋ]�E�P�E��P3��}�-Q���P�=�  ����t� ��u�E�j PSVW�i�����^�M�_3�[��R����U���0�H�3ŉE��ESW�}j[S�M�Q�M�Q�p�0�n�  ����u�g�����V������   V�u��u�L�����;������   �E�H3Ƀ}�-�E�������9;�t��+��M�Q�uPS��  ����t� �S�E�H9E������|+;E}&��t
�C��u��C��u�E�jP�uVW��������u�E�jP�u�uVW�Q�����^�M�_3�[��Q����U��j �u�   YY]�U���W�u�M��O���U�}��
��t���   � � :�tB�
��u��B��t4�	<et<EtB���u�V��J�:0t����   ��:uJ�BF���u�^�}� _t�E��`p���U��j �u�u�u�   ��]�U��QQ�} �u�ut�E�P� �  �M�E���E��A��EP�s�  �M�E�����U��j �u�   YY]�U����M�V�u�3N���u�P������e�F�P蘉����Yu��P�ǧ��Y��xu���E�����   � � �F���ȊF��u�^8E�t�E��`p���U��E�������Az3�@]�3�]�U��W�}��tV�uV�Qw��@P�>VP��D����^_]�Vh   h   3�V�z�  ����u^�VVVVV������V3������8���������(r�^�U��E��u裙���    �������]Ë@]�jh�u�(����u���u�A����  �m���� 	   �   ��xy;5��sq��������������D8��tSV�-�  Y�e� ����D8tV�U   Y�������� 	   ����}��E������
   ���)�u�}�V肨  Y�謘���  �ؘ��� 	   �������������U��VW�}W�h�  Y���tP����u	���   u��u�@Dtj�=�  j���4�  YY;�tW�(�  YP� ���u
�L����3�W脦  Y������������D9 ��tV����Y����3�_^]�U��V�u�F�t �Ft�v�!c���f����3�Y��F�F^]�jh�u�����}���u����� 	   �   ����   ;=����   �����E��߃�������D��ttW薣  Y3��u��E�����Dt(W�0�  YP�����u�L����u��t�*����0�W���� 	   ����u��E������
   ���!�}�u�W�ʦ  Y��(���� 	   �������� ����jh�u�����u���u�ǖ���  ����� 	   �   ����   ;5����   ��������������D8��tcV諢  Y�e� ����D8t�u�uV�_   �����腖��� 	   �F����  ����}��E������
   ���)�u�}�V��  Y������  �F���� 	   �1�����������U���  請  �H�3ŉE��E�M3�W����@�����D�����<�����,���9Uu3���  ��u试��!8�ܕ���    ���������  SV������������0������������\$�����t��u+�E�Шu�S���!8耕���    �k����L  ��@����D tjRRP��  ����@�����  Y���  ��0�������D��   �����@l3�9��   �����P��0���������4��@����������  9�@���t����  �����D���!�$����ʉ������4���9}�~  3���8���ǅ���
   ����  �	3���
����@�����0�������|8 t�D4�E�j�E�M��d8 P�Z��P�hn  Y��tD��D�����4���+�E����  jR��<���P�/�  �������  ��4���@��8����&j��4�����<���P� �  �������  ��4���3�QQ@��8���j��4����E�Pj��<���PQ������@���������k  j ��$���QP�E�P��0�������4�������  ��8���������,���9�$����!  ��@��� ��   j ��$���Pj�E�P��0����E�����4�������  ��$�����   ��,���G�   ��t��u3�3�f;������<�����8���������4�����8�����@�����t��uU��<����أ  Yf;�<����  ����@��� t$jXP��<���诣  Yf;�<�����  G��,�����8�����4���;E������#��0�������G�D4����D8   ��@����  ��@����  ��0�������D��U  ��D���3���8�������   ��<���9u��  3�+�<�����H�����@���;EsD�
B@��#�����
��@�����<���u��,����CA��#������<���CA��@������  r��������H���+�j ��(���PS��H���P��0�������4�������  �(�����D���9�(�����  ��<���+�;E��<����5����  �ʀ���   ��@���9u��  ǅ���
   ����� ��,�����+������H���;Es>�1������@���f;����ujYf���@���������f�3�������  r��������H���+�j ��(���PS��H���P��0�����,�������4�����8�����<�������  �(�����D�����<���9�(�����  ��@�����+�;E� ����  �]��$�������  ǅ���
   ����� ��$���+ʋ������H���;�s;�>������$���f;����uj^f�0��$�������f�8�������  r�3�VVhU  ������Q��H���+��+���P��PVh��  �@���8�����<�����4�������   3ɉ�@���j +���(���RP������������P��0�������4�����t��@����(�����4�����@���;����L���@�������4�����8���;�Q��$�����D�����+���<���;�������7j ��(���Q�u��D����4�����t
��(���3���L�����D�����uc��t$j[;�u�r���� 	   �3�����?V�<���Y�6��0������������D@t	�:u3�� �2����    �����  ����+�,�����^[�M�3�_�]D����U��W�}��u������    �������   �G����   �@��   �t�� �G��   ���G�  u	W�  Y��G��w�wW�����YP���  ���G����   �����   �G�uQW�����Y���t0W����Y���t$VW������W��������Y����Y^�����@$�<�u�O    �   u�Gt�G   u�G   ��O�A���������	G�g ���_]�jdhv����j�"k��Y3ۉ]�j@j _W����YY�ȉM܅�uj��E�PhH��S  ������U  ���=��   ;�s1f�A 
�	��Y�a$��A$$�A$f�A%

�Y8�Y4��@�Mܡ��ƍE�P���f�}� �)  �E����  ��M���E���E�   ;�|�ȉM�3�F�u�9��} j@W�\���YY�ȉM܅���   ����M���}ԋE؋U�;���   �2���tX���tS� �tM�uV����U���t8����������4���u܋��E؊ �Fh�  �FP�l��F�U��M�G�}ԋE�@�E؃��U�놉��=�����   ;�s$f�A 
�	��Y�a$�f�A%

�Y8�Y4��@�M���F�uЋM������]ԃ���   ����5��u܃>�t�>�t�F��F�   �F���uj�X�
�C�������P��������tE��tAW�����t6�>%�   ��u�F@���u	�F�Fh�  �FP�l��F�"�F@�F���������t
���@����C�<����E������   3��.����j��i��Y�VW���>��t7��   ;�s"���� tW�0����@��   �G�;�r��6�U���& Y�����|�_^�jh(v聿��3��u������u�ȉ���    ����������,V��S��Y�e� V�2   Y���}��ډ]��E������   �ǋ��p���Ëu�]�}�V�T��Y�U��$  ��~  �H�3ŉE�S�]VWS����3���Y������9{}�{jWWV�  ��������������;�|;�s
�����9  �����΋4�������������D$����C  ������������������u�C�������������+��������  �;��+s�C��  �������D  ����������������|
0 �������   ��{ ��  ���������������j �t,�t(S��  �������������������������������;|(�����;T,�����j ������Rh   ������R�4� ��������������������j WQS�V  ����������������������;��������������t3���N;�s*�<u�B�;�s�A�8
u���������A��uэ�����+�3��������������}  ����������������D�������t�K��9
uFA;�r����u��3��>  �C�u��
����    ������C�	  �{ u3���   ������+{���������{�D���������������   jj j �������,  ��������������������;�u$9�����u�C�8��8
uG@;�r��C    �_j RQ��������  �����4������,����   ;�w�Ct�C   ��t�{����������������������D������tG������u��+ǃ� ������������u��3��������M�_^3�[�<����U��V�uWV����Y�N�����u誅��� 	   �N ����  ��@t莅��� "   ��S3���t�^��t}�F�����N�F�����F�^�  u*�rO���� ;�t�fO����@;�uW���  Y��uV�
  Y�F  tz�V��B��F+�H�M�F��~QRW����������G�� �N�h���t���t�ϋǃ������������A tjSSW�A   #����t%�N�E��3�@P�E�EPW��������;]t	�N �����E[_^]�jhHv��������u؉u܋}���u�%����  �Q���� 	   �   ����   ;=����   �����E�߃�������D��tpW��  Y�e� �E����Dt�u�u�uW�g   ��������؃��� 	   虃���  �މu؉]��E������   ���+�}�]܋u�W�>�  Y��h����  蔃��� 	   �����֋��k����U��QQV�uWV�!�  ���Y;�u�b���� 	   �ǋ��D�u�M�Q�u�uP����u�L�P����Y�Ӌ�����������d0��E��U�_^��U���u����u�L��3���tP�ɂ��Y���]�3�]�U��V�uW�9EuI�}j�P;Mu+�y��YY���u3��.�E�    �6�u�7�9�����Q��y������tՉ�&3�@_^]�U��S�]��P�q����Y��u��߃�[]�U��M�Ix
��@��	Q�=���Y�Ћ�]�U����  �H�3ŉE��M�E��4��� �� ��� SW�}�����3ۍ�|�����p�����\�����P���ǅ(���^  ��`�����u�ف���    �ĺ������h  ��t��@@VurP����Y�Ⱦ�����t���t�у�����������B$u&���t���t��������������A$�t�\����    �G��������  �u�������4���3�3Ɉ�y�����l�����d�����8�������  �������T����������D�����P�cp��Y��tPN��d�����p�����d���VP�  YY���t	VP�I��YYG�P�*p��Y��u�d�����\�����l�����  �j%Y:��B  8O�/  ��\���3ɉ�<�����3�����L�����@�������[�����Z�����z�����j�����{������,�����F���H�����P�Eo������H���Ytf��@���k�
������z�����{�����tĈ�k�����`�����\�����l�����t������  ��������������������H�����   ��N��   t���*ty��Ft���It��L��   ��끊F<6u#�N�94u����,�����D��� ��T��� �W���<3u�N�92u���D���<d�<���<itx<o�0���<x�(���<Xu'������z�������z���������ht;��lt��wt��������F�8lu���w����Ǌ�{�������{�����z����������{��������㊍{����ქH��� ��\���2���x�����u�<Stƅ{����<Cuƅ{����:�� ��nt[��ct&��{t!��p�����d���P�#  ��d���Y��l������p���F��l�����d���������؉�`���Y�����  ��\�����@�����t�����t���g  ��o��  ��  ��c��  ��d�x  ��  ��g~*��it��n��  ��z��� ���  �Q  jd_�  3���-u��P���F����+u*��l�����p���I��t���G�6����؋�@���Y��`������l�����u	�����t�����P�l��Y��t�����tj��I��t�����t]��P�����L������4���P��|���P��P���P��(���PFV�?��������r  ��p���G��������P��`����l��Y닋�������   � � ��[���:���   ��I��t�������   ��p���G�Y�����P����؊�[������4���P��|���P��P���P��(���PFV��`�������������
  ��P�k���n��t�����I��t�����t`��P�����L������4���P��|���P��P���P��(���PFV�D��������w
  ��p���G��������P��`����k��YY��u���L��� �c  ��et	��E�U  ��t�����I��t������>  ��P����e��4���P��|���P��P���P��(���PFV����������	  ��p���G� �����Y��`�����-u9��P������4���P��|���P��P���P��(���PFV�f���������	  ���+u0��t�����I��t�����u��t������p���G������Y��`�����P�j���n��t�����I��t�����t`��P�����L������4���P��|���P��P���P��(���PFV����������	  ��p���G�=�������P��`����i��YY��u�O��l�����d������t��p���S�B��YY��L��� ��  ��z��� ��  ��P�����8��������Q��H���P� ��k���QHP�5���<��Ѓ��  ��uAǅ@���   ��t�����{�����~ƅj�����l�����H���I��l�����d������t��p���S��A��YY��l�����@��� t��t�����J��t�������  ��p���A��l�����d���������Y��`�������q  ��ctF��su��	|	���Y  �� u.��{�K  3ҋ˃�����B���L���[���3ȅ��&  ��z��� �  ��j��� ��  ��P��$����S  Y��t%��l�����p���@��l�����d����u���Y��%��������P�����ǅ ���?   �pt��$���P�� ���P趈  ��H���f�� �����f�����H���������ǃ�p��  ���s���HH��  ���  ��t1�;���  ��y����Ȁ�z��� ��  �����������  ��{�����~ƅj���B��\����:^uB��\���ƅ[����j �E�j P�4����\������:]u	�]B�E� �~��3����vB��\���<-uP��tL�
��]tEB��\���:�s����Ċ�����у�����D����̰;�|�փ�������D�2���Ȋ��у������D܋�\����<]u�����  ��\����W�����@�����-u	ƅZ������+u8I��t���u��t
���x����!��p���F��l�����d���������Y��`�����0��  ��p���F��l�����d����m�����Y��`�����xtb��Xt]ǅL���   ��xt&��@��� t��t���H��t���u��x���jo_�G  N��l�����d������t��p���S�>��YYj0[�  ��p���F��l�����d����������@��� ��Y��`���t��t�������t�����}��x���jx늋�H����@��H����E���F�?�����l���H��l�����d������t��p���S�>��YY��H���;��%  ��z��� �=  ��8�����c�.  ��j��� t
3�f��  �  �  ƅk�����@�����-u	ƅZ������+u2I��t���u��t��'��p���F��l�����d��������Y�؉�`�����x�����,��� �\  ���#  ��xta��pt\��P�)d��Y����   ��ou$��8��   ��T�����D�������T������g��T���j j
Q��D���Q�M����ȉ�T����F��P�yd��Y����   ��D�����T�������S��T�����D���������Y��D�����`�����L����CЙȋ�T����@��� ��D�����T���t��t���tR��p���F��l�����d����������Y��`��������N��l�����d������t��p���S�><��YY��D�����T�����Z��� �	  �ك� �؉�D�����T�����   ����   ��xt;��pt6��P��b��Y����   ��ou��8��   ��<������5��<���k�
�*��P�Cc��Y��td��<���S������؋�<���Y��`�����L������Ã�@��� ��<���t��t���tL��p���F��l�����d����������Y��`����N���N��l�����d������t��p���S�3;��YY��<�����Z��� t�؉�<�����F���#�L����)  ��z��� uE��8�����<�����,��� t��H�����D������T����H���k����ɋ�H���t��f���y�����\�����l�����G��y�����\����m:�u8OuG��p���F��l�����d�����������GY��`�����\���;�ul��P�+L  Y��t&��p�������Y�G��\���;�u(��l�����d������u�?%uA�nu;���������/��p������t	VP��9��YY���tV����t��p���S��9��YY��4���u��P����<��Y��8������;�u��u8�y���t������� t
������ap�^�M�_3�[�'����U��SV�u�u��������Y���t��Q�`��Y��u�^��[]�U����V�   V�g��Y�M�A��t	�I�q��I�A�A�A   �A�a �^]�jhhv�v���3��}�j�O��Y!}�j^�u�;5�}S������tD�@�tP�/��Y���tG�}��|)������ P�0����4��~;��Y���$� F��E������   ���7���Ë}�j��O��Y�U���$�M��u��#���E��t�M��ESVW��t�}��t��|��$~�p���    ������  �}�3ۉ]��p�t~�E�P��jP�)  �}܃�����   ���H����t�F�ʋE�]���-u����M�F���+t�M��}�]�E����C  ���:  ��$�1  ��u��0tj
_�0�<xt<Xtj��j_�
��u��0u�<xt<Xu	�N�M������3����E�E܉U����   �U��E����H�ȃ�t	�E���0�%  tD�M��A�<��w�� ���;�s-�M��;�ru;E�v�E����t���؊�E�M�F랋EN�U��U���u��t�u3��I������u��u:��t��   �w��u';�v#�mn���U�� "   ��t����j ��[��ߋE��t�0��t����E��t�M�3ۀ}� t�M�ap�_^��[��U��=� j �u�u�uuhx��j ������]���3Ʌ�������Ã%� �����������U���SQ�E���E��EU�u�M�m��Y�  VW��_^��]�MU���   u�   Q�7�  ]Y[�� jh�v�����5��<���t�e� ���3�@Ëe��E������   �jh�v����譴���@x��t�e� ���3�@Ëe��E������k���腴���@|��t������h���8����U��V�u��������E  �V\W�}��99t�����   ;�r�   ;�s99t3Ʌ��  �Q���  ��u�a 3�@��   ��u�����   �ES�^`�F`�y��   j$_�F\���d� ���   |�9�  ��~du�Fd�   �   �9�  �u	�Fd�   �u�9�  �u	�Fd�   �d�9�  �u	�Fd�   �S�9�  �u	�Fd�   �B�9�  �u	�Fd�   �1�9�  �u	�Fd�   � �9� �u	�Fd�   ��9� �u�Fd�   �vdj��Y�~d�	�q�a ��Y�^`���[�3�_^]�U��csm�9Eu�uP����YY]�3�]�U��QQ�=�� u�j���SVWh  � �3�WS�$����5��=����t8u���E�P�E�PSSV�[   �]��������?sE�M����s=��;�r6R�a����Y��t)�E�P�E�P��PWV�   �E���H����=��3�����_^[��U��ES�]V�# �u�    �EW�}��t�8���E3ɉM�>"u3�����F�ȉM�"�5���t��G��E��PF�k��Y��t���t��GF�E��t�M��u�< t<	u���t�G� �N�e �> ��   �< t<	uF��> ��   �U��t�:���U�E� 3�B3��FA�>\t��>"u3��u�} t�F�8"u���3�3�9E���E���I��t�\G���u���tA9Mu< t8<	t4��t*��P�<j��Y��t��t��GF���G���tF��F�o�����t� G��-����U_^[��t�" �E� ]Ã=�� u�B���V�5�W3���u����   <=tGV�_F��FY����u�GjP�\_����YY�=����tʋ5�S�> t>V�*F���>=Y�Xt"jS�+_��YY���t@VSP�T������uH���> uȋ5�V�3���%� �' ���   3�Y[_^��5���3���%�� �����3�PPPPP�n����U����H��e� �e� VW�N�@��  ��;�t��t	�УL��f�E�P�h��E�3E�E��`�1E���1E��E�P���M�3M�E�3M�3�;�u�O�@����u��G  ��ȉH��щL�_^��U��QW����3���tuV��f9t��f9u���f9u�SPPP+�P��FVWPP�@��E���t7P�#^����Y��t*3�PP�u�SVWPP�@���u	S�p2��Y3�W� ����	W� �3�[^_��VW�Ti�Ti����t�Ѓ�;�r�_^�VW�\i�\i����t�Ѓ�;�r�_^�U���5(��<���t�u��Y��t3�@]�3�]�U��E�(�]�U���(3��E��E�90�t�5���<�����ީ�E��   V;���  ��  ���  ��   jZ+���   H��   ����   H��   ����   HtN��	�#  �E�   �E�PB�E�u� �E�]�� �E��]�P��]���Y����  �f��� "   ��  �E�LB�E�u� �E�]��E�   � �E��]�P��]���Y�  �E�   �E�LB��E�DB�V  �U��E�DB�l����E�@B�;  �U��E�@B�Q����E�PB놃�tfHtWHtHHt/���  ��	t���8  �E�TB��   �E�\B��   �E�PB�E�u� ���   �E�PB��   �E�   �������E���   �E�   �E�dB�����������   �$����E�@B��E�DB��E�LB��E�lB��E�tB�u����E�|B�i����E܄B�]����E܌B�E�u� �M��� �E�]�� �]��.�EܐB���EܔB���EܘB�E�u� �E�]�� �]���E��]�P�E�   ��Y��u�/d��� !   �E��^�Ë�8�A�J�S�\�h���t�������������j
��  �|�3��U��QQSV���  V�5 ��;  �EYY�M�ظ�  #�QQ�$f;�uT�3  YY��~-��~��u#�ESQQ�$j�6  ���qVS�W;  �EYY�c�ES��������\$�$jj�?�(  �U��E��������DzV��S���;  �E�YY��� u�S�Ƀ��\$�$jj�3  ��^[��U���  �H�3ŉE��ESV�uW�}�u������3��؍������������������������������������������������������������1���b������������������
  �@@ucP�����Y�ȃ��t���t�у������������B$��
  ���t���t���������������A$��b
  ���Z
  �3��Љ��������������������������������������
  ������������@����������	  �A�<Xw�����B���3���������ǸB��������������������������	  �$�}3���������؉������������������������������������L	  ���� tF��t9��t/HHt���������-	  ���������	  ���������	  �����ˀ   ������*u/�������������������  ���؉�������������  ������k�
�����������������ȉ������  3��������  ��*u+������������������������r  ��������f  ������k�
�����Љ������>  ��ItE��ht8��������lt��w�,  ��   ������8lu@��   �������������� ������������ <6u�������4u�ǃ��� �  ����<3u�������2u�ǃ����������<d��  <i��  <o��  <u��  <x��  <X��  3��������3�������������P��P�19  YY��t8������P�������������  ���������A���������������b  ������P�������������  ����  ����d��  �Q  ��S��   t|��AtHHtVHHtHH�  �� ǅ����   ��������������@�   ���������������������2  ǅ����   �  ��0  ��   ��   �������   ��0  u��   �������������������t�ʋ7����������  �S  ��u�5�ǅ����   �ƅ�t3�If9t����u�+����<  ��X��  HHtp���'���HH�$  ����������  t0�G�Ph   ������P������P��z  ����tǅ����   ��G�������ǅ����   ��������  �����������t3�p��t,� ��   t�+���ǅ����   �  3ɉ������}  �5�V�i:��Y�k  ��p��  ��  ��e�Y  ��g�K�����itd��nt%��o�=  ǅ����   ��y[��   �������M�����������x  ���   �������� tf���ǅ����   �z  ��@������ǅ����
   �� �  u��   ��  �����������3��  u��guVǅ����   �J;�~������=�   ~7��]  W��R��Y��������������t
���������
ǅ�����   ����������������G�������������P��������������������P������������VP�5���<��Ћ�����   t!������ u������PV�5���<���YY������gu��u������PV�5���<���YY�>-�(�����   ������F����ǅ����   j���s�����HH��������k  j'X������ǅ����   ���|���Qƅ����0������ǅ����   �^�����3��������� t��@t�G���G����@t
�G���ȋ���O�����@t;�|;�s����߁�   �������� �  u����������y3�B�����   ������;�~�Ћ��u�������u��J�����������t=�������RPWQ�/t  ��0����������������9~������������������N밋������E�+�F��������   t6��t�>0t-N�������0�!��u�5����I�8 t@��u�+Ɖ����������� ��  ��@t5��   t	ƅ����-���t	ƅ����+���tƅ���� ǅ����   ������+�����������+���u������P������Wj �   ��������������������Q������P������P�  ����t��u������P������Wj0�  �������� ������t}��~y��H�������Pj�E�P��������P��������u  ����u?9�����t7������������P�������E�������P�r  ����������������u��(����������#������������Q������PV�8  ����������x#��t������P������Wj ��   ����������������tP�#��3�Y������������������������������������������� _^[t
�������ap��M�3��	�����W���    蚐������ɋ�� ����-�������$U��U�B@t�z t-�Jx��M������ERP����YY���u�E��]ËE� ]�U��V�u��~W�}W�uN�u�������?�t���_^]�U��V�uW�}��G@�Et� u
�M�E�N�& S�]��~@�EP�EW� PK�K����E���E�8�u�>*uPWj?�/����E����˃> u�E�[_^]ø�ø�ø�ø���U��M��u�lV���    �W���jX]á��3�]�U��M��u�BV���    �-���jX]á��3�]�U��M��u�V���    ����jX]á��3�]�U����E�e� V��u��U��j^�0�Ҏ������  j$h�   P�~���E����t�S��@�E���
|��@W��rjY;�|���&A�v�U��j^�0���  Wj h�3�PS�{	  ��F�E��p�+  ���  ���M�jd_�u�j��}�h�����ȋƙ��+ȋƙ�������������E�������RP�b��+�j h�Q �RP�b���u���3�G��E|��s?�M�À3����� %  �yH���@u
����}��u��l  ��}���u9�ÀQ �� �+�M���%  �yH���@u
����}��u��l  ��}���u�}��}j h�Q VS�O�  j��G�h����RP��a����}� �8�u���W3�@9Q}@9�|�H�G+��Ej h�Q �W�p�0�*  j��Y���j h  VS�W�  j��G�h����RP�~a���j j<�VS��  �g  �Gk�<+؉3�_[^��jh�v�n����=<� u,j�2��Y�e� �=<� u�K  �<��E������   �y����j�83��Y�jh�v����j�1��Y�e� �u�&   Y���u��E������   ���6���Ëu�j��2��Y�U��QS�E�3�P�]�����Y����  9]��m  V�uW�N3�G;��u;���&  9@���   ���P���P���P���Pf9��u���SP���P���PQW����P���SSPQSW�h  �����,P���P���P���Pf9��u���SP���P���P�vW����P���SSP�vSS�  ��,�NjXjZ3�jC_��k}jXj
_3�jB[j j j jj j RPQjj��  3�PPPjPPSW�vjP�  ��X�=������V;�};�|$;� ;�~ ;�}3�@_^[��;�|�;��;�~;�}3���Nk�<N3�k�<i��  ;�u;������;�����SSSSS�a����j0hw����3ۉ]̉]ԉ]�]܉]؉]�j�/��Y�]������E��E�P�����Y����   �E�P����Y����   �E�P����Y����   �1A���Eȉ@���������hTC�n  Y���}���tx8tt�8���tPW�O��YY��t(�8���tP���YW��-��@P�,G��YY�8���u�E�   �   WW�-��Y@P�58�����������   SSSSS�O����8���tP�L��Y�8�hH��$�3�F�����   �5@��H�k�<�M�f�=�� t���k�<ȉM�f�=�� t�����t�u�+��k�<�E���]܉]؍E�PSj?�E��0j�hL�S�u��@���t�}� u
�E�� �X?��E�� ��E�PSj?�E��pj�h��S�u��@���t�}� u�E��@�X?��E��@��uԋu�������0�u������0�u������0�E������a   �}� ��   jWj@�u��6�.  ������������?-u�E�   GW����Y��i�  �M�<+t<0|<9G��3ۋÉE̋}�j�s.��YÀ?:uBGW���Yk�<�M�ȉM��<9G�<0}��?:uGW���Y�M�ȉM��<9G�<0}��}� t�ىM�? t �E�   jWj@�v��-  ����t������]܋F��u������0�u������0�����U����e� �}S�]VW����   %  �yH���@jd�E���  Yu	�Ù����u��l  �����t�E���� ���E����4��E��+  ���Gj���C������i�m  ��%���+��C�����������^���M��k�+�;U���E�����   �}� u��jd�Y����u��l  ���  ����t�E����	�E��8�;�~I+��E%  �yH���@u��jd�Y����u��l  ���  ����t�E�<� ��
�E�<�4�} �E$k�<E(k�<E,i��  E0�}u�=��������_^[�ã���E�P�=���F���Y��uF�E����i��  ȉ��y�� \&����� \&;�|+�����������j j j j j �C����V�Ɠ������u�+L���    3�^Ã~D uj$�B��Y�FD��t܋FD^��������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� ������SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ��������������U���0���S�ٽ\�����= � t��  ��8����   [����ݕz������U���U���0���S�ٽ\����= � t�#  ��8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8����3  �   [�À�8�����=� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �xC�����������hC����s4��C�,ǅr���   �pC�����������`C����v��CVW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�Rf  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����K   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[��������̀zuf��\���������?�f�?f��^���٭^�����C�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����C�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����C���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-�C��p��� ƅp���
��
�t���U��E�����]�U����M�S�u�����]�C=   w�E苀�   �X�n�����E�M���QP��  YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�E�PQ�E�P�E�jP�  ����u8E�t�E��`p�3���E�#E�}� t�M��ap�[��U��Q�e� V�E�P�u�u��  ������u9E�t�WE����t
�NE���M����^��U��V�u��t�U��t�M��u3�f��!E��j^�0�~����^]�W��+��f��If��tJu�3�_��u�f���D��j"��U��Q�H�3ŉE��MSVW3���u�E� �@�E��3�9E WW�u���u��   PQ�D��؅�u3��   ~A�����w9�]   =   w辍�����t����  �P������Y��t����  �������t��PWV�� ����SV�u�uj�u�D���t�uPV�u�H���V����Y�Ǎe�_^[�M�3��Q�����U����u�M������u �E��u�u�u�u�uP��������}� t�M��ap���U��} u�u���Y]�V�u��u�u���Y3��MS�0��uFV�uj �5��(��؅�u^9,�t@V�e���Y��t���v�V�U���Y�QC���    3�[^]��@C�����L�P�EC��Y����(C�����L�P�-C��Y�����U��V�uW3���tj�3�X��;Es��B���    3��<�uS�]��t	S�Cx��Y��VS������YY��t;�s+�V�j P�j�������[_^]�U��V�u��tj�3�X��;Es�B���    3��Q�u��uF3Ƀ��wVj�5��d��ȅ�u*�=,� tV�N���Y��uЋE��t�봋E��t�    ��^]�U��E��VW�}3���t���?  3�f�S�]��u�B���    ��z������  �u�M��}����E����   9��   u(9u��   �f��< ��   F��;ur���   �u���WVSj	�p�D�����   �L���zuR�M���*I�M����t'�E�P��P�A  Y���EYt@�8 t%�M�@�E��u��u+�WP�E�Sj�p�D���u!�+A��� *   3�f��99��   uS�V��Y���&VV���VSj	�p�D���u��@��� *   ��p��}� t�M�ap���[_^��U���S�]VW�}3���u��t���u�@��j^�0�y���   3�f��E��t�0�u�M�������9]w�E=���v	�o@��j�C�M�QP�uW�-��������u��t3�f��G@���0�:@��t,;�v!�}�t3�f��*@��j"^�0�y���jP��^3�f�LG��M��t��}� t�M��ap�_��^[��U��j �u�u�u�u�u������]�U���,�H�3ŉE��ES�]VW�}3��E�}�u���t��u3��   ��u�?���    �x������  �u�M������M�Eԅ���  9��   u4����  ��   f9�T  ��1f���f���v  F;�r��l  �xtua��t"�ǋ�f90t��Ju���tf90u��+���C�EԍU�RVSQSWV�p�@�������   �}� ��   �E�|0� �  N�  �U�RVSQj�WV�p�@�����t9u���   �w���   9u���   �L���z��   ����   �E�M�Q�M�V�qt�U�RjPV�q�@��Ѕ���   9u���   ����   ����   �:;���   �ƉE��~�M�D�9����   �E�@G�E�;�|�E���E�;�r��j��=��� *   ����&9��   u"�f��t��   f;�w2��F�f��u���0�M�QVVVj�WV�p�@���t
9u�u�x���=��� *   ����}� t�M܃ap��ǋM�_^3�[�������U��QV�u3�W�}�E���t.��t.��t�S�]��t���9}w�E=���v �3=��j�Y��t��&=��j^�0�v�����k�uP�uV�4��������u��t� ��<��� �E@��t5;�v'�}�t� ;�w��<��j"^�0��u�����jP��Y��M��D0� ��M���t���[_^��jh(w�Cr��3ۋ�u�j����Y�]����}�;=���   ������tV�@�uF�@ �  u=�G���w�GP�$��Y��t~���4�W���YY�����@�tPW����YYG떋��u��Mj8�2��Y�ȡ�����t7h�  ������ P�l������� P�(����4��u�^��t�f �  �^�^��^�N��E������   ���q��Ëu�j�E��Y�U��QQS3�!U�V�u3�W�=p��E��F�> t��<at-<rt"<wt�[;���    �Ft��3��+  �  �3ۃ���	  ��3�AF�����  �E   ���  ����S��   tv�� ��   ��tRHtC��t-��
t��u�9E���   �E�   ���   �ˀ   �   ��@��   ��@�   �E�   �   ��u���������π   �t�}� uh�E�   �� �b��TtP��t;Ht+��t�������� �  u9�� @  �7��u-B�������*��u B�� @  ��� �  u�� �  ��E��t3���F���������E�����   �F�> t�jVh�C��Y  ���������j ��X�F8t��>=�r���F8t�jh�CV��Z  ����u����   �Cjh�CV��Z  ����u����   �$jh�CV�Z  ������������   �F�> t��> �����h�  �u�ES�uP�)Y  ������������E3ɉH��H�H�M�x�H_^[�����������������SVW�T$�D$�L$URPQQh�'d�5    �H�3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�RT  �   �C�dT  �d�    ��_^[ËL$�A   �   t3�D$�H3�����U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�S  3�3�3�3�3���U��SVWj RhF(Q蚗  _^[]�U�l$RQ�t$������]� U��   �1-  �H�3ŉE�S�]��������u�7���    �yp������  VS�����3�Y������9C}�CjPV��  �ȃ���������y�����  ��������������ƃ����������T$����C  ������u
+K���  �3W��+{�C�������z  ���  ����������������|0 ��������   ��{ u���>  ���������������j �t,�t(S�����������������������;t(��  ;T,��  j ������Rh   ������R�4� ����m  j ������S��  �����T  ������;��F  ��������t3���O;�s*�<u�B�;�s�A�8
u���������A��uэ�����+��1�U  ����������������D�������t*�K������;΋�����s�������8
uG@;�r���������u���   �C�u��c5���    �   �C��   �{ u3���   +ss����������������D���������   jj �������   ��������;�u�C�0��8
uF@;�r��C    �Uj Q�������r   ����y����W�   ;�w�Ct�C   ��t�s����������������D������tF��������u��+΀�u��_^�M�3�[������jhHw��i���u���u�4���  �>4��� 	   �   ����   ;5����   ��������������D8��tcV��?  Y�e� ����D8t�u�uV�_   �������3��� 	   �3���  ����}��E������
   ���)�u�}�V�;C  Y��e3���  �3��� 	   �|l������ii���U��V�uV�"B  Y���u�e3��� 	   ����LSW�u3�W�uP�,��؃��u�L�����tW�3��Y����������������d0���_[^]��5���<��U��E���������� �]�j$hhw�|h��3ۉ]�3��}؋u��Pt��jY+�t"+�t+�t^+�uH�8z�����}؅�u����d  �E�������^�w\V�S  YY���E� �V�ƃ�t6��t#Ht�`2���    �Kk����E��������E��������E� �� �3�C�]�P�<��E܃���   ��uj�e����tj �J��Y�e� ��t
��t��u�G`�EЃg` ��uA�Gd�E��Gd�   ��u/��A�щUԡ�A�;�}&��k��G\�d B�Uԋ�A��j �8��M��E������   ��u �wdV�U�Y��u�]��}؅�tj ���Y�V�U�Y��t
��t��u�EЉG`��u�ẺGd3��g���U��M��AV�u9qt��k�E��;�r�k�U;�s	9qu���3�^]�U���EW��������Dz	��3��   Vf�u�Ʃ�  u|�M�U���� u��tj�ٿ�������Au3�@�3��EuɉM��y���M�O�Et�f�u�U���  f#�f�u��t� �  f�f�u�Ej QQ�$�1   ���#j ��QQ�$�   �������  �����  ^�E�8_]�U��QQ�M�E�E�]����  ��%�  �f�M��E���U��}  ��Eu��u@]Á}  ��u	��ujX]�f�M��  f#�f;�uj���  f;�u�E�� u��tj��3�]�U��E� tj��t3�@]ètj��tjX]������]�S��QQ�����U�k�l$���   �H�3ŉE�V�s V�CP�s�   ����u&�e��P�CP�CP�s�C �sP�E�P�  �s ���s�c����= � Yu)��t%�CV���\$���\$�C�$�sP�  ��$�P�V  �$��  V�  �CYY�M�3�^�������]��[�U���S�]V�����t�Etj�  Y����  ��t�Etj�n  Y����u  ����   �E��   j�K  �EY�   #�tT=   t7=   t;�ub��M����Ю��{L�H��M�����{,�Ю�2��M�����z�Ю���M�����z���������������   ����   �E��   W3���tG�M���������D��   ��EPQQ�$�����E�U��� ������E=����}3���G�W��3�����AuB�E�����f�E��E����;�})+ȋE��E�t��uG���E��E�t   ��E��m�Iu��E��t���E��3�G��_tj��  Y�����t�E tj ��  Y���3���^��[��U��= � u%�u�E���T$���\$�$�uj�W  ��$]��,��h��  �u� !   �]  �EYY]�U��j �u�u�u�u�u�u�   ��]�U��E3ɉH�ES�H�E3ۉH�MCW��t�E��  �	X��}��t�E��  ��H��t�E��  ��H��t�E��  ��H��t�E��  ��H�MV�u�����3A��1A��M���3A��1A��M����3A��1A��M����3A��1A��M����3A#�1A��  ����t�M�I��t�E�H��t�E�H��t�E�H�� t�E	X��   #�t5=   t"=   t;�u)�E��!�M���������M��������E� ���   #�t =   t;�u"�E� ���M�������M�������E�M��3���� 1�E	X �}  t,�E�` �E� �E�X�E	X`�E�]�``�E��XP�:�M�A �����A �E� �E�X�E	X`�M�]�A`�����A`��E�XP�  �EPjj W�T��M�At�&��At�&��At�&��At�&��At�&ߋ��������� t/HtHtHu(�   � �%����   ���%����   ��!������� tHtHu!��#�   �	�#�   ��}  ^t�AP���AP�_[]�U��E��t�����w�T)��� "   ]��G)��� !   ]�U��U�� 3ɋ�9��t@��|������M��tU�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E��   �E�P�r������uV�Y���Y�E�^��h��  �u(�   �u�=����E ����jh�w�;^���=ľ|[�E�@tJ�=� tA�e� �U�.�E� �8  �t�8  �t3��3�@Ëe�%� �e��U�E������
�࿉E�U�^���U��Q�}����E���U��Q��}��M�E#E��f#M�f����E�m�E���U��QQ�M��t
�-Я�]���t����-Я�]�������t
�-ܯ�]����t	�������؛�� t���]����U��Q��}��E���U��=� uu�U��u�w'���    �b`������]ËM��t�SVWjA_jZ+�[�
f;�rf;�w�� ������f;�rf;�w�� ����f��tf;�t�����_^+�[]�j �u�u�   ��]�U����M�SV�u�����]��t�u��u��&���    ��_�������   �E�W���    uBjAYjZ+�Z�3f;�rf;�w�� ������f;�rf;�w�� ����f��t:f;�t��3��M�QP��R  ����M�QP�[��R  �����vf��tf;�t�����+�_�}� ^[t�M��ap�����U����u�M������E��M���   �H% �  �}� t�M��ap���U��j �u����YY]�U��3ҋ�9Ev�Mf9t	@��;Er�]����U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�?C  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ���D�   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z���D������������D�����   s���D���D������������D�����   v���D�U��VW�}��t�M��t�U��u3�f��#��j^�0�\����_^]Ë�f�> t��Iu��t�+��f��Rf��tIu�3���u�f��f#��j"�U��U�MV��u��u9Mu&3��3��t�E��t��u3�f���u��u3�f�� #��j^�0�\����^]�SW�ً����u+��f�3�vf��t%Ou�� +��f��[f��tOtJu��u3�f���_[�{������u�E3�jPf�TA�X�3�f��"��j"�U��E��x!��~��u���������]��t"���    �_[�����]�U���$�H�3ŉE��ES�8�VW�E�E3�W�E��Ӌ��u�����E�9=���   h   Wh�D�4�����u$�L���W�h  h�D�8������S  h�DV������?  P��h�DV�����P��hEV�����P��hEV�����P�ӣ���th8EV���P�ӣ��u�����t�E��tP�0�9}�tjX�   9}�t�5��<�j����<�;�tO95�tGP���5��E��ӋM�E��t/��t+�х�t�M�Qj�M�QjP�U��t�E�u�u��    �0��;�t$P�Ӆ�t�Ћ���t��;�tP�Ӆ�tW�Ћ��u�5��Ӆ�tV�u��u�W���3��M�_^3�[�������U��U�MV��u��u9Mu!3��.��t�E��t��u���u��u� �E ��j^�0�1Y����^]�SW�ً����u+ފ�3F��tOu��+��C��tOtJu���u���_[u����u�EjP�D� X�� ����j"�U��QQ�H�3ŉE��ES� V�@W3�VV�u�E��u�3J���؃���u3��   ~Ej�3�X���r9�]   =   w��h������t����  �P�������Y��t����  �������t�SW�u�u��I������t VV9uuVV��u�uj�WV�u��@���W����Y�ƍe�_^[�M�3��[�����U����u�M������u�E��u�u�uP�������}� t�M��ap�������U��ES�H<�V�A�Y��3��W��t�}�p;�r	�H�;�r
B��(;�r�3�_^[]��������������U��j�h�wh �d�    P��SVW�H�1E�3�P�E�d�    �e��E�    h   �|   ����tT�E-   Ph   �R�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE� 3Ɂ8  �����Ëe��E�����3��M�d�    Y_^[��]�������U��E�MZ  f9t3�]ËH<�3��9PE  u�  f9Q��]�U��E� �]Ã%x� �U��V�u����   �F;D�tP�f���Y�F;H�tP�T���Y�F;L�tP�B���Y�F;P�tP�0���Y�F;T�tP����Y�F ;X�tP����Y�F$;\�tP�����Y�F8;p�tP�����Y�F<;t�tP�����Y�F@;x�tP�����Y�FD;|�tP����Y�FH;��tP����Y�FL;��tP����Y^]�U���S�]3�VW�M��]�M�9��   u9��   u���M��8��  jPj�����YY�u��u3�@�K  j������Y�}���u	V�!���Y�ރ' ���    �y  j���Y�E���uV�����W�����Y�σ  ���   �FPjW�E�jP�J���M��QjW���E�jP�J����E��PjW�E�jP�J����E��PjW�E�jP�vJ����E��P��PjW�E�E�jP�YJ����E�� PjPW�E�jP�BJ����E��$PjQW�E�jP�+J����E��(PjWj �E�P�J����E��P��)PjW�E�j P��I����E��*PjTW�E�j P��I����E��+PjUW�E�j P��I����E��,PjVW�E�j P�I����E��P��-PjWW�E�j P�I����E��.PjRW�E�j P�I����E��/PjSW�E�j P�mI����E��8PjWj�E�P�VI����E��P��<PjW�E�jP�<I����E��@PjW�E�jP�%I����E��DPjW�E�jP�I����E��HPjPW�E�jP��H����E��P��LPjQW�E�jP��H�����t)�]S�a���S������E�P������E�P������������U���<0|<9,0�B�: u��"<;u��F��v�> u���}jY�8�󥋃�   �u� ����   �}��@�F���   3ɋ@�F���   A�@0�F0���   �@4�F4�E����t����   ��tP�$��{x t"�sx�$���u���   �����sx����YY�E��Cx���   ���   3�_^[��U��V�u��tY�;8�tP�����Y�F;<�tP����Y�F;@�tP����Y�F0;h�tP����Y�F4;l�tP����Y^]�U���S�]3�VW�]�E�9��   u9��   u���E��8��D  3�FjPV�u����YY�E��u���n  ���   jY��j����Y�E���u�u����3�Y@�A  3��89��   �K  j�|��Y�E����   �u�8���   jW�E�jP�F���M��QjW���E�jP�F����E��PjW�E��E�jP�|F����E��0PjW�E�jP�eF����E��P��4PjW�E�jP�KF�����t%�u�n����M��Y�u�I����M�Q�@����E�YY�w�U����<0|o<9k,0�B�: u�}�u�M�3�@���t��{| t	�s|�$��{x t"�sx�$���u�sx��������   �����YY�E��Cx�{|���   3�_^[��<;u���F��v�> u�녡8��u��<��F�@��F�h��F0�l��F4�a���U��V�u���n  �v�b����v�Z����v�R����v�J����v�B����v�:����6�3����v �+����v$�#����v(�����v,�����v0�����v4�����v������v8������v<�������@�v@������vD������vH������vL������vP������vT�����vX�����v\�����v`�����vd�����vh�����vl�����vp�����vt�x����vx�p����v|�h�����@���   �Z������   �O������   �D������   �9������   �.������   �#������   �������   �������   �������   ��������   ��������   ��������   ��������   ��������   ��������   ������@���   �������   �������   �������   �������   �{������   �p������   �e������   �Z������   �O������   �D������   �9������   �.������   �#������   ������   ������  ������@��  �������  �������  �������  �������  �������  ������   ������$  ������(  ������,  ������0  ������4  �{�����8  �p�����<  �e�����@  �Z�����D  �O�����@��H  �A�����L  �6�����P  �+�����T  � �����X  ������\  �
�����`  �������^]�U��SVW�}���    t?3�hd  CS�	����YY��u���KWV�I   YY��tV�A���V����YY�߉��   ��X����   =X�t�   P�$����   3�_^[]�U��QQSV�uW�}���   ��u�����  S�\���e� ��`  �GPj1S�E�jP�u��A���OQj2S���E�jP�
A����GPj3S�E�jP��@����@��GPj4S�E�jP��@����GPj5S�E�jP��@����GPj6S�E�jP�@��Wj7S��E�jP�@����P��G Pj*S�E�jP�@����G$Pj+S�E�jP�{@����G(Pj,S�E�jP�g@����G,Pj-S�E�jP�S@����P��G0Pj.S�E�jP�<@����G4Pj/S�E�jP�(@����GPj0S�E�jP�@����G8PjDS�E�jP� @����P��G<PjES�E�jP��?����G@PjFS�E�jP��?����GDPjGS�E�jP��?����GHPjHS�E�jP�?����P��GLPjIS�E�jP�?����GPPjJS�E�jP�?����GTPjKS�E�jP�n?����GXPjLS�E�jP�Z?����P��G\PjMS�E�jP�C?����G`PjNS�E�jP�/?����GdPjOS�E�jP�?����GhPj8S�E�jP�?����P��GlPj9S�E�jP��>����GpPj:S�E�jP��>����GtPj;S�E�jP��>����GxPj<S�E�jP�>����P��G|Pj=S�E�jP�>������   Pj>S�E�jP�>������   Pj?S�E�jP�o>������   Pj@Sj�E�P�X>����P����   PjAS�E�jP�>>������   PjBS�E�jP�'>������   PjCS�E�jP�>������   Pj(S�E�jP��=����P����   Pj)S�E�jP��=������   PjS�E�jP��=������   Pj S�E�jP�=������   Ph  S�E�jP�=����P����   Ph	  S�E�j P�z=������   Pj1S�E�jP�c=������   Pj2S�E�jP�L=������   Pj3S�E�jP�5=����P����   Pj4S�E�jP�=������   Pj5S�E�jP�=������   Pj6S�E�jP��<������   Pj7S�E�jP��<����P����   Pj*S�E�jP�<������   Pj+S�E�jP�<������   Pj,S�E�jP�<������   Pj-S�E�jP�w<����P����   Pj.S�E�jP�]<������   Pj/S�E�jP�F<������   Pj0S�E�jP�/<������   PjDS�E�jP�<����P����   PjES�E�jP��;������   PjFS�E�jP��;������   PjGS�E�jP��;������   PjHS�E�jP�;����P���   PjIS�E�jP�;�����  PjJS�E�jP�;�����  PjKS�E�jP�q;�����  PjLS�E�jP�Z;����P���  PjMS�E�jP�@;�����  PjNS�E�jP�);�����  PjOSj�E�P�;�����  Pj8S�E�jP��:����P���   Pj9S�E�jP��:�����$  Pj:S�E�jP��:�����(  Pj;S�E�jP�:�����,  Pj<S�E�jP�:����P���0  Pj=S�E�jP�:�����4  Pj>S�E�jP�k:�����8  Pj?S�E�jP�T:�����<  Pj@S�E�jP�=:����P���@  PjAS�E�jP�#:�����D  PjBS�E�jP�:�����H  PjCS�E�jP��9�����L  Pj(S�E�jP��9����P���P  Pj)S�E�jP��9�����T  PjS�E�jP�9�����X  Pj S�E�jP�9�����\  Ph  S�E�jP�|9����P�_^[��Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ��U��UV�uW�:�+�u+�f��t���:�+�t�_^��y����~3�A��]�U��Q�MS3�VW��f9t3�}���f��t��M��M��f;U�t���f��u�3҃�f9u�_+�^��[��U��E��u]ËM�UVHt�2f��tf;1u��������	+�^]�U��ES�VWf��t*�}���f��t��f;�t���f��u����f��u�3�_^[]�U���   �H�3ŉE�V�u��P����N  jUP�4��YY��~*��P���P��	��@P��P���P��P  jUP��������u�M�3�^�5�����3�PPPPP��A���U��V�u�6�	���v�����@�F�r	�������@�~ YY�FtjX��6�~   Yj jh7X�F�|2�����F   t�F   t�Fu�f ^]�U��V�u�6�	�������@Y�FtjX��6�"   Yj jhUZ�F� 2�����Fu�f ^]�U��M3҅�u3�]����f��Arf��Zv	���f��wB���]�U���   �H�3ŉE�SV�u��x����8O�����   j@�K��ɍ�|��������P��  QV�2������u	!C@�g  W��|���P�s�����YY��������   j@��|���P�C���#�  PV��1��������   ��|���P�3����YY��u*�K  V����@PV��P  jUP��������tF�/  �Cu;�{ t�s��|���P�3��1  ����u�K��CuV�L  Y��t�K뜋C�   #�;���   �K���h�   ��|���#�P��  QV�1������u	�c 3�@�[��|���P�3�����YY��u<�K   3�9{tJ�K   f9�P  uV���@PV��P  jUP���������u\�C���Ѓ�_�M�^3�[�g����� 9{t��3����Y;Cu�V�y  Y��u��3������3�����YY;�t���x����x���3�WWWWW��>���U����   �H�3ŉE�VW�}� M�����   jx�N��ɍ���������P��  QW� 0������u!F@�A�����P�6�����YY��u"W���@PW��P  jUP���������u�N�F���Ѓ��M�_3�^�x����� 3�PPPPP�>���U��V�u��tWf�> tQh�RV����YY��t@h�RV����YY��u&j�EP�EP  h   P�I/������t/�E^]�V�b3  Y��j�EP�EP  h  P�/������u3��ЋE��u�^]�%��U����H�3ŉE�V�uj	�E�PjYV��.������tj	�E�VP���������@�M�3�^芺����U��V�u3�WB3���xPS��tJ�M�7�+�����k��E�4�E�0�n�����YY��u�E�M��ȋE��
y�s���{;�~�[3���_��^]�U��QSVW�5K���]���   3ɍ�P  �E�f����   �~�N��f9tWjh P�O�����3ɋVf9tF�f9t����������~ Yu2Vj@hPE��������t�3�Vf9t�g���������������Y3�9~�  ��   VP�������YY����   ����  ��   ����  ��   ��P�������   �E��t�0�}����   �u���   3�f��v��@P�u�jUS�G���������   j@Wh  S�-������tnj@���   S��   h  P��,������tMj_S�!1  YY��uj.S�1  YY��tj@S��   jP�,������tj
j��   PV�/  ��3�@�3�_^[��3�PPPPP�;���U����   �H�3ŉE�SV�uW�aI�����ZI�����  V�  Y���   ��ɋ�h�   ����������P��  QV�����u!@�6�����P���   �����YY��uV�  Y��t	��w�w����Ѓ��M�_^3�[谷���� U��V��H�������   �������Y�j@h^���   ����E^� u�  ]�U��VW�H�����   �6�����v�����@�F����}�����@�F�g �~ YYtjX��6�   Yjh`�F����   t�   t�u�' _^]�U��V�H�������   �F�������@Y���   tjX����   �"   Yjh�a���   ����E^� u�  ]�U��M3����f��Arf��Zv	���f��wB���]�U����   �H�3ŉE�SV�uW�sG�����   �hG�����  V�  Y�K��ɋ�h�   ����������P��  QV�����u�' 3�@�t  �����P�s����YY����   h�   �����P�C���%���  PV�����t������P�3�����YY��u�  �w�R�uP�{ t0�s�����P�3�*  ����u��w�3�����Y;Cu�w����uV�  Y��t����w��   #�;���   �K���h�   ����������P��  QV���������������P�3����YY��u"�   9CuF9CtA�3�J���Y;Cu4Wj�"�{ u8�{ t2�����P�3�����YY��uWPV�  ����t�   � u�w����Ѓ��M�_^3�[�}����� U����   �H�3ŉE�SV�uW�E�����   �uE�����  V�   Y�K��ɋ�h�   ����������P��  QV�����u!@�`�����P�3�!���YY��u
9Cu4Wj�"�{ u2�{ t,�����P�3�����YY��uWPV�'  ����t	��w�w����Ѓ��M�_^3�[褳���� U��UV�
3�f��t9Wj_�A��Rf;�w����  ��A�f;�w����  �Ƀ������
f��u�_��^]�U��V�u��tRf�> tLh�RV����YY��t;h�RV����YY��u!j�EP�Eh   �p�����t*�E^]�V�Q+  Y��j�EP�Eh  �p�����u3��ՋE��u�^]�%��U��M3�f;��Rt����r�3�@]�3�]�U��QVW�C���uj���E�P�΁��  h   ��   Q�����u3��,;u�t$�} t���   ��������   ������YY;�t�3�@_^��U����H�3ŉE��ESV�u�E�EW�E��:C�����   3�jP�E�P�d������C���M����  ��u�M�  �   ���   �{3ɉ3���tf9t��RWHPh P�.�����3ɉM����tgf9tb���tf9t�E�P�#����	�E�P�����}� Yup��RSHPhPE���������tM���t3�f9t�E�P�������E�P�T�������tf9t�E�P����Y��E�  ����E�E��}� ��   �E�P��   ���#�V������YY����   ����  ��   ����  ��   ��P�������   j�u������t�E��t�0jU��P  P�u��#���]����tVjU��   P�u��k#���=����j@Sh  �u��ׅ�t0j@���   Ph  �u��ׅ�tj
j��   QV�y'  ��3�@�3��M�_^3�[�$����������U��W�=ľ��   �}ww�U�����fn��p� ۹   #σ����+�3��of��ft�ft�f��#�uf��#���ǅ�EЃ������Sf��#���3�+�#�I#�[��ǅ�D�_���U��t93���   t�;�Dǅ�t G��   u�fn�f:cG�@�L�B�u�_�ø����#�f��ft �   #Ϻ������f��#�uf��ft@��f����t����뽋}3�������ك��E���8t3�����_��U��UV�uW�z��u�|���j^�0�h1�����   �} v�M� ��~���3�@9Ew	�J���j"��S�^�0�Å�~���t��G�j0Z�@I���U�  ��x�?5|�� 0H�89t�� �>1u�B�S�<���@PSV�Ӣ����3�[_^]�U���(�H�3ŉE�SV�uW�u�}�M��X����E�P3�SSSSV�E�P�E�P��1  �E�E�WP�	'  �ȋE��(�u��t��uj�
�u��tj[�}� t�M��ap��M�_^��3�[謭����U���(�H�3ŉE�SV�uW�u�}�M��̪���E�P3�SSSSV�E�P�E�P�j1  �E�E�WP��+  �ȋE��(�u��t��uj�
�u��tj[�}� t�M��ap��M�_^��3�[� �����U��QQ�ES�PVW�x� �������  �� �  ����� �   ��}��E���t���  t�� <  �%��  �!��u��u�E!P!f�x�X��<  3����M���������]���E�s���x&�������������  �y�}�}��E�s�f�{_^[��U���0�H�3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���uЋ���f��7  �u܉C�E��E��C�E�P�uV�2�����$��u�M�_�s^��3�[�۫����3�PPPPP�.������������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��U��M�E������#�V�u�����t$��tj j �z@  YY��9���j^�0�%-�����Q�u��t	�V@  ���M@  YY3�^]�j��&��Y�jh�w�)���}����������4���~ u0j
�#���Y�e� �~ uh�  �FP�l��F�E������*   ��������������P�(�3�@�q)��Ë}j
�-���Y�jh�w�)������u�e� j�2���Y��u��j  j����Y�e� 3ۉ]؃�@�B  �<������   �}����   ;���   �GuW� u0j
�K���Y�E�   � uh�  �GP�l��G�e� �/   �E܅�u�GP�(��Gt!�GP�,���@뇋u�]؋}�j
�P���YËE܅�u��G����+4����������u���uC�+���j@j ����YY�ȉM���te������ ���   ;�sf�A 
�	��a ��@�M��ۋ����u�����΃�������DV�����Y��u����u��E������   ����'��Ëu�j����Y�U��EVW��x`;��sX��������������Dt=�<�t7�=X�u3�+�tHtHuQj��Qj��Qj��<������3���c���� 	   �$����  ���_^]�U��M���u�
����  �6���� 	   �B��x&;��s������������Dt�]�������  ������ 	   ��)�����]�U��MSW��x\;��sT��������������<�u:�=X�V�uu�� tItIuVj��Vj��Vj��<�����43�^��z���� 	   �;����  ���_[]�U��M��������������P�,�]�U��M���u�/���� 	   �8��x$;��s������������D��@]������� 	   ��(��3�]�U���SV�u��t�]��t�> u�E��t3�f�3�^[��W�u�M��K����E����    u�M��t�f�3�G�   �E�P�P�a���YY��t@�}��t~';_t|%3�9E��P�u�wtVj	�w�D��}���u;_tr.�~ t(�t�13�9E��3�GP�u�E�WVj	�p�D���u�������� *   �}� t�M��ap���_�6���U��j �u�u�u�������]�U��Q������u
�>  ������u���  ��j �M�Qj�MQP�@���t�f�E��jhx�9$���u���u�R����  �~���� 	   ��   ����   ;5����   ��������������D8����   ����;E�@u������  �#����    �vV����Y�e� ����D8t�u�uV�_   ����������� 	   �����  ����}��E������
   ���)�u�}�V�U���Y������  ����� 	   �&������#���U���(�ESV�uWj�Y3��}��M�u�;�u�=����8�j���� 	   �O  ���0  ;���$  �����؋�������M�D�]ܨ��  �����v������8�����    ��  ����  ���  9}u	����!8�ҊD$����E��HtHu���Шtۃ���E�E��d���Шt����sj^V�K���Y�E���u�����    �]����    �v  jj j �u��h���M������D(�E��T,�M����M��DH�E���   �T��
t|��tx�3��P���GN�} �U��D
tZ����D%<
tK��tG����BjN�}�U�_�D%
u+����D&<
t��tj_����j
BY�U�N�L&�u�y������E�Ytq����D�tc�E�P�4����E���tL�}uFj �E�P�E�����V�u��4�D���u�L�P�8���Y����E��  �E� �M��8�E���j �M�QV�u��4� �����  �M����  ;���  �U���4���D���W  �}�m  ��t�M��9
u�$��D�E����8�E��M�;��  jY���<��   :�t	�FG�   �E�H;�s�G�8
uj
X����   �F���xj �E�Pj�E�P���G�4� ���u
�L���u|�}� tv�U����DHt#j
Xj8E�u�F�&�����E�F�D�;u�uj
X8E�u�FjY;}��D����Kjj�j��u�lf���U��j
X8E�t�jY�F�ыU�jY�F�Ƌ���D�@u�D���F�E���+��}�  ����   N���xF�   ��3�B��� u�]���;�rNB���� t�]�������u�I���� *   �����@;�u��\�E����DHt7�F�D�E��|�����D%�E�F��u�����D&F+���ڋjRP�u�]e�����E؋}���P�u+�VWj h��  �D������M����E�3ɋ��;�����L0�E��]�;EtP蜳��Y���t�����n  �}� ty�u��Ǚ+������΍G;�sUj�E   _�f;Et3f;�tf�������B�;�sj
��Xf9tjXP_f���;�r���E����L�E���+�����d�����t�M�j
Zf9�U�u�$��D�E����8�E؉M�;��_  jY�E   ���f;E�&  f;�tf��'�E����;�s(j
Zf9W�U�uj
X��f���   f������   j �E�Pj�E�P������4� ���u�L�����   �}� ��   �U����DHtRj
Xjf9E�uf����3Xf�����E��D����E��D%���j
Y���L&jY;}������l;u�uj
Xf9E�uf�����jj�j��u�4c���U��j
Xf9E�t�jYf���뷋U�jYf���멋���D�@u�D�	f�f����E���+�������L�j^;�u�M���� 	   �����0�������m�����3������3��������8����� 	   ������_^[����������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� �����������U��SVWUj j h�z�u�E  ]_^[��]ËL$�A   �   t2�D$�H�3��m���U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�zd�5    �H�3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�zu�Q�R9Qu�   �SQ���SQ���L$�K�C�kUQPXY]Y[� ���U��QQ�E���]��E��ËH���3�9l����U���S�]W�}��u��t�E��t�  3���E��t��V�����v�����j^�0����X�u�M��B����E�3�9��   u`f�E��   f;�v9��t��tWVS�4������v���� *   �k����0�}� t�M��ap���^_[�Å�t��t_��E��t��    �ӍMQVWSj�MQV�u�p�@��ȅ�t9uu��E��t����L���zu���t��tWVS觟���������j"^�0�����q���U��j �u�u�u�u�������]�U��=�� V�5��u3��cW��u95��tS�2  ��uJ�5����t@�} t:�u�����Y���'Q赿��Y;�v��<8=uW�uP��2  ����t�����u�3�_^]Ë@���S��QQ�����U�k�l$���   �H�3ŉE��CV�s��W��|���Ht+Ht$HtHtHtHHtHuzj��   �nj�
j�j�j_Q�FPW�)�������uG�K��t��t��t�e����E��F����]����E��FP�FPQW��|���P�E�P�
�������|���h��  Q�L����>YYt�= � uV�+��Y��u�6�ڷ��Y�M�_3�^茗����]��[�jh0x�����e� 3��u������u����j^�0�������^��3�9E����tރ} t�E%������@tɃe� �u�u�u�u�uV�E�P�U   �����}��E������   ��t�������Ëu�}��}� t%��t�������������d��6����Y�U��Q�e� �E�P�u�3��YY��u�����V�u �u�u�u�u��u�u��  �u����9����� ��^��U��j�u�u�u�u�u�������]�U��j �u�u�u�   ��]�U���V�u��u3���   SW�u�M��`����E�3�9PuV�u�u�7��������   �]��t�}��u�����    ��������   ��U�N��C�Dj �]�Zt4��u��]����Dum����I���u�������f�C�ɉ]���U���G�Dj Zt��u����N��t�����f���Gf;�uf��t�]����q����҃�J�}� _[t�M�ap���^��U��j �u�u�u�   ��]�U����M�SVW�u�A����}3҅���  �M�9QuW�u�u��/  �����i  �u��t�]��u�j����    �U�������A  ��E�E���OF�D�u�tl��u��U��D�  ���f����   ���u�U��X�e��f	E�E��F�u�f���E�f;qrf;qwfq�/f;qr)f;qw#fq�f�u����Dt��  �E�f�u���E��E��C�DtI��u�U�b�O��t��e���f	E��E���C�Ef;Arf;AwfA�8f;Ar2f;Aw,fA�&f�E��j �D
�UZt�E��  �Ef�Ef;�uf��t�u���������҃�J�}� _^[t�M��ap�����U���V�������t"h$Zh����P�������u����\�u��������Et2�e� �e� �E�E �E�E�E�E�P�u�E�   �u�u�u���E j P�u�u�u�u�u��^��U���8S3��E�W�]��]��E�   �]�t	�]��E��
�E�   �]��E�P�_0  Y���  �M� �  ��u�� @ u9E�t�M�������   �+�tHHt*Ht#�������E�������j[��������  ��� ��t��   t���U���   @��   ��}��EVj^jZ�U�+�t6+�t)+�t +�t��@uu��   ����E���E�   ��U���E�   ��]��%   �   ;�(t!��t=   t=   tJ=   u"���Fj�j^�==   t3=   t(=   t%�������E������j[�������  j��3�F��   �ÉU�E���   t�����#E����x3�B�U���@t��   �M��   �E��}���   t	��   �U���    t   �E��� t   �
��t   �E�������}����u!�)�������S����    �H���� ^_[���u��E�u��    V�E�P�u��u��u�������E���us�M��   ���#�;�u1�Et+�u��E��u�����VP�u�M�Q�u��������E���u2�������������d��L�P����Y������q  P�����uB�������������d��L���V�N���Y�u�� ���u��\����    맃�u�M�@�	��u�M��u��7�O����U�YY���������������T�������������U��d$��M��$H�E���   ����  ����   jj�j��7�MU����#ʃ��EԉU���u�����8�   tS�7��?�������j�E�P�7�]����������uf�}�u�u��u��7��*  �����t�SSS�7��T��#����t��U��M���  �� @ u�E�% @ u�� @  �ȉM��% @ = @  tD=   t)= @ t"=   t)= @ t"=   t= @ u�E����%  =  u	�E���]���   ��  �]���@��  �E��   �#�=   @��   =   �t[;��l  ���d  jY;��  ��v���  �F  QSS�7��S�������   SSS�7��S��#���������j�E�P�7���������������M�jZ;�t����   ��﻿ u	�E���   ����  ����  u�7�3>��Y�����j[��  ����  uJSSR�7�VS��#���������E��   ����   jY;�v6���"���QSS�7�S�����tSSS�7�S��#����uQ�����jY�E���HtHu=�E���  �jY�E�﻿ �M؋�+�P�E��P�7�1?�������������M��;�ً������������D$2E�$0D$�7�M��������������D2$��$
ȈL2$�M8]�u!��t�������������L �M�u��   ���#�;�u}��tx�u�� ��u��E��u�����jP�u�V�u���������u2�L�P�L����������������d��7�y���Y�����������������
�������SSSSS�%���U��Q�=� W��   �}3�����   �U��u������    ���������t�M��t�SVjA[jZ^+щu��jZ^�
f;�rf;�w�� ������f;�rf;E�w�� ����Ot
f��tf;�t�����^+�[�j �u�u�u�   ��_��U���SV3�W9u��   �]��u�J����    �5�������   �}��t��u�M�輇���E�9��   uQ�MjAZjZ^+߉u��jZ^�;f;�rf;�w�� ������f;�rf;E�w�� ����ItDf��t?f;�t��8�E�P�P�G   ���E�P�P�7   ���M���[�t
f��tf;�t�����+��}� t�M�ap���_^[��U����  ��f9E��   V�u�M������u싆�   ��u�M�A�f��wf�� ������   jf9Us*�u�W   YY��u	�E����M���   �����M�Qj�MQRP���������u	�E����E��}� ^t�M�ap���U��Qf�E���  f;�u3��ù   f;�s�ȡ$��H��E�Pj�EPj�H����#E����M#���U��}
�Eu
��yjj
�j �u�u�uP�   ]�U��MV��u�6���j^�0�"������   �} SWw����j^�   �U3���f���@9Ew	�����j"�ދEj"���^;�w�3��ҋU�E��tj-Xf�3�@�y�E�ڋM�ߋ�3��u�U�ЋE��	v��W���0f���A��t;Mr�;M�Mr3�f������0�t
����� 3�f����f�f�f�����;�r�3�_[^]� U��j
j �u�C(  ��]�S��QQ�����U�k�l$��Kf�S�� �=ľ|H��fn��p� fp� ��%�  =�  w>�of��fu�fu�f��f����u4����f;�t���f��u�3�f9��H#��"�f;�tf��t������E����3������]��[�U���D�H�3ŉE��MS�A
��% �  �E��A�E��A�E�����  V���?  W�}��3ۉ}��U��E������u%���9\��u@��|��  3��}𫫫j[�  �t��u��}�H��H�U܉E̋��j�^#�����]ԉUā�  �yI���A+�3�@����j����u�^�D����   �����ЅD���9\��u
B;�|��   �E̙jY#�ЋE���%  �yH���@+�3�@��j��]�_�EȋD���M�ȉM�;ȋE؋�r;E�s3�A�M�J�D��x.��t'�D���ˍx;��]ԉ}؋�r��s3�A�M�J�D��yՃ���MЋUċ���!D���B;�}�}��΍<�+�3�����M�9]�tA�p���+t�;�}3��}𫫫������;��  +U܍u�UЋ�}�������EċEХ%  �yH���@�EЃ���ǋ}Ћ���j �]��ЉE�X+�j�E�^�T����#E؋���M���U�C�T��E�;�|ߋE����U�j+ЋE�3�Y���;�|��D���E���\����Iy�M�A���������Uԁ�  �yI���AjX+��EЋM�3�@���D����   �����ЅD���9\��uB;�|��v�}̋ǙjY#������  �yO���G�D��+�3�G��j��ˉ}���}�;��E�_r;E�s3�AJ�D��x(��t!�D���ˍx;��}���r��s3�AJ�D��yۃ���MЋUԋ���!D��B;�}�}��΍<�+�3�����x�A���������E؁�  �yI���A�M����j �]��]�Y+��׉ẺM܋T������M�#�U��T���M����E��E�@�E�;�|׋u؋����U�j+�Y3�;�|��D����\����Iy������;l���   �x�3��}𫫫�M�   ����������É�  �yI���A�����j X+��M��׉]��E؋T������M�#���U��MȉT��C�E�;�|ߋű����U�j+�Y3�;�|��D����\����Iy�5��5l�3�C�   �5���e�����x����������uȉE؁�  �yI���A��j �]���X��+ÉM��׉E܋T������M�#���U�F�T��E���|ߋ}؋uȋ����U�j+�Y3�;�|��D����\����Iy�}�jX+x��ȋE������%   ��|�u���@u
�E�w���� u�7�M�_^��3�[�v�����U���D�H�3ŉE��MS�A
��% �  �E��A�E��A�E�����  V���?  W�}��3ۉ}��U��E������u%���9\��u@��|��  3��}𫫫j[�  ����u��}�H��H�U܉E̋��j�^#�����]ԉUā�  �yI���A+�3�@����j����u�^�D����   �����ЅD���9\��u
B;�|��   �E̙jY#�ЋE���%  �yH���@+�3�@��j��]�_�EȋD���M�ȉM�;ȋE؋�r;E�s3�A�M�J�D��x.��t'�D���ˍx;��]ԉ}؋�r��s3�A�M�J�D��yՃ���MЋUċ���!D���B;�}�}��΍<�+�3�����M�9]�tA�����+��;�}3��}𫫫������;��  +U܍u�UЋ�}�������EċEХ%  �yH���@�EЃ���ǋ}Ћ���j �]��ЉE�X+�j�E�^�T����#E؋���M���U�C�T��E�;�|ߋE����U�j+ЋE�3�Y���;�|��D���E���\����Iy�M�A���������Uԁ�  �yI���AjX+��EЋM�3�@���D����   �����ЅD���9\��uB;�|��v�}̋ǙjY#������  �yO���G�D��+�3�G��j��ˉ}���}�;��E�_r;E�s3�AJ�D��x(��t!�D���ˍx;��}���r��s3�AJ�D��yۃ���MЋUԋ���!D��B;�}�}��΍<�+�3�������A���������E؁�  �yI���A�M����j �]��]�Y+��׉ẺM܋T������M�#�U��T���M����E��E�@�E�;�|׋u؋����U�j+�Y3�;�|��D����\����Iy������;����   ���3��}𫫫�M�   ����������É�  �yI���A�����j X+��M��׉]��E؋T������M�#���U��MȉT��C�E�;�|ߋű����U�j+�Y3�;�|��D����\����Iy�5��5��3�C�   �5���e����������������uȉE؁�  �yI���A��j �]���X��+ÉM��׉E܋T������M�#���U�F�T��E���|ߋ}؋uȋ����U�j+�Y3�;�|��D����\����Iy�}�jX+���ȋE������%   �𡔱u���@u
�E�w���� u�7�M�_^��3�[�|����U���|�H�3ŉE��E�E��E�E�3�S3�@V�E���W�}��]��]��]��]��]���]�9E$u�g����    �R���3���  �M�щU���� t��	t
��
t��uA��A���{  �$����B�<wjXI���E$� ���   � :ujX����+tHHt����  3�@�j� �  X�U��jX�]��3�@�E��B�<v��E$� ���   � :uj묀�+t+��-t&��0t���C�3  ��E~��d���"  j�|���Ij�t����B�<�P����E$� ���   � :�R�����0�c����M���  3�@�E���0|*�E��u���9��s	��0@�G�F�A��0}�u��E���E$� ���   � :�I�����+�t�����-�k����E���3�@�E��E��E���u��0u�E��HA��0t��E��E���0|%�u���9��s��0@�GN�A��0}�u��E����+������-������C~��E�������d�������I�  3�@��0�E���	����j�/����A��E��B�<wj	������+t"HHt�������j����j���X�U������j����3�@�E���A��0t���1����   몍B�<v���0�9] t"�A��E���+t�HH�q����M��jX�}���j
XI��
�p����A3�@�E������9,k�
������P  
�A��0}���Q  ���9�A��0}�I�E��U��
�M�����  ��v�E�<|���E��M�OjAX�M���M�����  O8u
HAO8t��M��M�QP�E�P�  �U�����y�ދE�u���uu�E���u+u��P  �,  �������  �����`����  y
� ��ރ�`9]��  3�f�M���  �΃�T���E��u�����  k�ȸ �  �M�f9r��}����M���M��M��y
�U΋�3�% �  �E���  #�#��]�����  �]ԉ]؉]܉u�f;��+  f;��"  ���  f;��  ��?  f;�w�]��  f��u$F�E�����u�u�}� u�}� u3�f�E���  f��uF�A����u�u	9Yu9t�j��_�E��U؉}��}���~\�uč4F�A�E���� �E���}����}�z��]�;z�r;}�s3�@��E��z���tf��E�����I�E�����M��}��E���@O�E��}�����u��U܋}ԁ��  �U�f��~;��x2�E؋ȋ����U��E���Ҹ��  ����}ԉU��U�f���f��i���  �f��y]�]��������E���E�tC�M؋����M��m�	E��E���������M��U܉E؉}�u�j �ۉU�[tf��3�Gf�f�Eԋ}��f�EԺ �  f;�w���� �� � u@�Eփ��u4�Eډ]փ��u f�E޹��  �]�f;�uf�U�F�f@f�E��@�EڋM��@�E֋M���  f;�sf�E�u�f�EċE؉EƉM�f�u��3�f9E���H%   � ���Ẻ]ĉ]ȋE��u����1����E��MċUƋu����23��ˋË�Ӎ_�#��  �   �j��ˋË����Ë�j�ˋ�[�}�E�f�f�G
�W�w�ËM�_^3�[�t���Ð��K���֛7���Ӝ6��x�m�B�U���   �H�3ŉE��US�]V� �  #��u3ɸ�  A#�W�]��E������E������E����?�U��E�f��t�C-��C �}f��u:����   9}��   3�f�� �  f;�����$ �C�Kf�C0 ����  f;���   �E�   �f��M;�u��t�   @uh�Z�Gf�}� t=   �u��u0h�Z�;�u%��u!h�Z�CjP��g��������  �C�h�Z�CjP�g��������  �C3��9  �֋�i�M  ����������Hk�M����ȋE�E�3��M���f�E��ٸ����`3�f�u�}�M��E�   �E���  �E��?  ���!  y�ٸ ���`�M����
  �u��U�u��}���T�E�����  k�ȸ �  ��x���f9r��}ĥ��Mĥ�MƉ�x����y
�E�}�1E�%�  ���  �E�Ǿ �  !u��}����E�N�]��]��]�]��}�f;��J  f9u��u��=  f;}��3  f;}�w�]��<  f��u G�E�����}�u��u��u3�f�E��$  f�}� uG�A����}�u	9Yu9t�j��^�E��U�u��u���~o�u��F�q�M��E���|����8����B��]��48;��u���r;�s3�F��u��B���tf��E���|�������I�E���|��������x����u��E���@N�E��u����w����}��E��u����  �E�f��~;��x2�E�������E�E��������  ���u��E��E�f���f��q���  �f��ye�]��������3҉}��}��E�B�U�tG�M�����M��m�	E��E���������M��]��E�u�u�j �]����}�[tf��f�f�E��u��f�E� �  f;�w���� �� � u@�E���u4�E��]���u f�E����  �]�f;�uf�M�G�f@f�E��@�E��M��@�E�M���  f;�s f�E�}�f�E��E�E�u��M�U�f�}��!3�f9E���H%   � ���E��Ӊu��U�u��E��M���������U�u��E�����?  f;���  �E��ȋEڋ�3��� �  �}���  #�#ωE������  �]��]��]�]��}�f;��@  �E�f;E��3  f;}��)  f;}�w�]��2  f��u G�E�����}�u��u��u3�f�E��  f��uG�E�����}�u�}� u�}� t���j�U��M�X����~X�}��E؍<W�E��}����ЋA��]��<;�r;�s3�@��E��y���tf��}��E�����N�}��E�����U��E���BH�U��E�����}��u����  f����   �]��]���x,�E�ȋ����E�������  ����]��u�f��Љ]��U�j [f��~[f�M� �  f;�w���� �� � ��   �E�����   �E��]�����   f�E����  �]�f;�u|� �  f�E�G�|�U���  �f��y���������}��}��E��E�tG�]�ˋ��������������M��]�U�u�j ���}��u�[�M���3�f��@f�f�M��U��<���f@f�E��@�E��u��@�E��  f;�s f�E�}�f�E��E�E�u�U�u�f�}��3�f9E���H%   � ���E����E�M��E��}f�t6���}���/3�f�� �  f9E�����$ �A3�@�A�A0�Y�  �}�jX;�~�E��}������?  3�j�}�f�E�]�_�ʋ���������Љu��]�Ou�}�j �]��U�u�[��y7�߁��   ~-�]��ʋ�������������O�]�u����]��U�u�3ۋu��E��~@�ω}��M��E�����   �u��}ĥ���}��ʋ����ЋE����4 ���ǋ������ЋE����8�M�;�r;�s�B��;�r��s3�A�ɋM���tF�Eȍ<;�r;�sF�U�u�ҋ����U��U��?Ћ����6��M��E���0��E�AH�U�M��]�E���~�E�E��>����u��}��A���<5|C�	�99u�0I;�s�;�sAf���E�*Ȁ��H�Ɉ\3�@�M�_^3�[�k���À90uI;�s�;�s΋M�3�f�� �  f9E�����$ �A3�@�A�0����3�SSSSS�x����U��M3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tƋѻ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t;�u �  ]Ã�@]�@�  ]�U�����}�f�E�3ɨtjY�t���t���t��� t���t��   SV���ֻ   W�   #�t&��   t��   t;�u��   �
����   ��   t;�u��   ���   ���   ��t��   �}�E����#�#��;���   V�=  ��Y�E��m���}��E�3��tj^�t���t���t��� t���t��   �Ћ�#�t*��   t��   t;�u��   ���   ���   ��   t��   u��   ���   �   ��t��   �=ľ��  ���]�E�3Ʉ�yjY�   t���   t���   t����t���   t��   �л `  #�t*��    t�� @  t;�u��   ���   ���   j@%@�  [+�t-�  t+�u��   ���   ���   ��#}��#��;���   P�$���P�E����YY�]�E3Ʉ�yjY�   t���   t���   t���   t���   t��   �п `  #�t*��    t�� @  t;�u��   ���   ���   %@�  +�t-�  t+�u��   ���   ���   ��3�Ω t��   ������_^[��U��M3���t@��t����t����t����t�� ��   t��V�Ѿ   W�   #�t#��   t;�t;�u   �   �   �с�   t��   u���_^��   t   ]á�����t���tP� ��3�PPjPjh   @h�Z������U��QV�5��W3��}��bWWWWj�PWW�@�����t`jW�#���YY�E���tOj j WPj��63�WW�@���t.�E�WP�  YY��y9}�t�u��z��Y�}������u�_^���u��z��Y�����U��j �u�u�u�   ��]�U����M�VW�u��b���E��u3��   �M��t�U��u�"����    ���������[����;�v�����    ������@�}� u�uPRQ��
  �����%�wPRPQh  ��  �E�P������� ��t�p��}� t�M��ap�_��^��U��=� VuH�} u芮���    �u��������>�} t����9uv�c����    �N������^]�  j �u�u�u�   ��^]�U����} ��   SVW�u�M��a���}������t�]��t�M;�v������    ������M�E����    uQSW�
  �����2+���M�QP�׹������M�QP�ȹ����C�Mt��t;�t�+��}� t�M��ap�_��^[��3���U���SVW�}3�jVVW�މu���)���ʉE�#����M���tYjVVW��)����#����tC�u�E+�E���   ����   h   j��P�d��E��u�����    ������ _^[��h �  W�?  Y�E��E�Y��|��   r�   ���P�u�W��������t�+��E�E�x#ȅ�t���j����8u蔬���    ���	]��u�W��   YY�u�j ��P�P��f��n|��shj �u�uW��(��#�����C���W����YP�������H��؋�#ȉE����u&�����    �٫�����L��#]���������j �u��u�W�j(��#���������3������U��M��u�ū���    ����jX]át��3�]�U��SV�u��������W�<���L7��%�   �E�D7$��ЋE��= @  tY= �  tI=   t*=   t#=   uP�ɀ�L7����D1$$��D1$�4�ɀ�L7����D1$$�����L7��ɀ�L7����d0$��} _^[u� �  ]���ҁ� �  �� @  ]�U��E�M����t���u�ª���    ����3��ËE��t
��|���$�SVW�93ۍq��>��jW�����YY��u�Ef��-u���f��+u�>���E��E��u6W�~  Y��t	�E
   �L�jxYf;�tjXYf;�t	�E   �0jX�E��u%W�C  Y��u�jxYf;�tjXYf;�u�~�����3��u�U�E�W�  ��Y���uHjAXf;�wf��Zv&j�G�Yf;�v�E��}���u_��t�u3��   jY�G���f;�w�� ��ɋM�E�;�sʋ}����E�;�ru;U�v�}���E���t������>���m����u�u@�ȃ�t��   �w��u-�����v%�4���� "   �E��t����j �[�Á������t�7�t��_^��[��U��j �u�u�u������]�U���S�]3�V�N@  W�E���S�S9U�@  �ʉM�U��U�U��}䥥��u��}������������ҋ��������E�������3ɉ�s�{�E;�r;E�s3�A���t��3ɍp;�r��s3�A�s��tG�{�U�3���M�;�r;�s3�@�K��tG�{�U}�u�e� ���������?��M҉�s�C�9�u��:�E�}�M;�r;�s3�B��U����t'�N3�;�r��s3�B��K�M�u���t@�E�C�C�EH�E�s�E��������N@  3�9Su.�S��������ЋE�������  ��E���tۉS�s�S�� �  u4�;�s���������E�������  ��E��� �  tى;�s�S_^f�C
[��U����E�e� W��u�����    ���������tS�V��t\j=S��  ��YY�u��tI;�tE�=��3�8F���E�;=��uW��  ���E�Y�=����ul9}t$9=��t������tL�w����    ���^[_�Å���  j�����Y�����t߃  �=�� uj�ߜ��Y�����t  �=����t���+�PS�  ��YY��xW�? tR�4��q���}� Yu���}�' �   �D���F�<� u�����?snjV�5�������}����tY����R�}� ��   ��y�ލF;��0���=���?�%���Pj�5��远�����������}�d� ���' 몋}�} tjjS袂��Y��P誛����YY��tPSS艂��Y��PV��O������uc��+�M��E�A�����#�PV�H���u�M������� *   V�p��Y�}� t
S� p���' Y�E��t���S��o���}Y�' 3��`���3�PPPPP������U��V�u3ɋƅ�tN9t	�@A�8 u�SW�AjP������YY�߅�uj	�k���Y���t+�P�>  ���Y�>��u�' _��[^]�U����V��W���t0�}WP�u���������u��<=t ��t�����uً��+�����_��^]�+5������U����M�SVW�u�W���E��u3��   �M��t�U��u�ѣ���    ���������h����;�v豣���    �����M�}����   ��u�u�VPRQ�T��������-�wPRPQh  �E�SP������ ��u�b����    ��p��}� t�M��ap�_��^[�����������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��U��f�Ej0Yf;���  f��:s��+�]ú�  f;��^  �`  f;��^  �J
f;�s��+�]ú�  f;��A  �J
f;�r�f	  f;��+  �J
f;�r͍Qvf;��  �J
f;�r��Qvf;��  �J
f;�r��Qvf;���   �J
f;�r��Qvf;���   �J
f;��y����f  f;���   �J
f;��_����Qvf;���   �J
f;��G����Qvf;���   �J
f;��/����P  f;�r{�J
f;������Qvf;�rg�J
f;�������Pf;�rS��Pf;�������@  f;�r=�J
f;��������  f;�r'�J
f;��������0f;�r��0���  f;���������]�U��} u3�]�SW�u�i~���xW�v����YY��t�uWS�K������u
���3�_[]�3�PPPPP������U��j �u�u�   ��]�U����M�VW�u�[T���U��u趠���    ����3��Z�}�3�9wu>�uR�
���YY���A���D8tB���t0�������9Mu�r����9Et	B�
f��u���9Eu��}� t�M��ap�_��^���%X��%�����̋T$�B�J�3��lV����l�yr������̋T$�B�J�3��LV���\m�Yr������̋T$�B�J�3��,V���m�9r������̋T$�B�J�3��V���n�r������̋T$�B�J�3���U����m��q������̋T$�B�J�3���U���dn��q������̋T$�B�J�3��U����i�q������̋T$�B�J�3��U����i�q������̋T$�B�J�3��lU���Tl�yq������̋T$�B�J�3��LU����k�Yq������̋T$�B�J�3��,U����j�9q������̋T$�B�J�3��U����k�q������̋T$�B�J�3���T���Dj��p������̋T$�B�J�3���T���Lk��p������̋T$�B�J�3��T����j�p������̋T$�B�J�3��T����o�p������̋T$�B�J�3��lT����o�yp���M��C?���T$�B�J�3��IT����p�Vp���T$�B�J�3��.T����s�;p���������h���<H��Y�����h ��,H��Y�����h��H��Y�������������h ���G��Yù ��%>��h����G��Y�h����G��Y�h����G��Y�h����G��Yù<���=��h���G��Y������@����������D����������H���������U��Q�=Դ uX�̴��t!����5ܴ�@<Q�@�Ѓ��̴    �ش��t#�٧���ش�E��E�P�H������ش    ��]ù ��=������@������\���?��?E���<��r=��                                                                     �y �y 
z z ,z � � hz |z �z �z �z �z �z �z { { 2{ H{ Z{ j{ v{ �{ �{ �{ �{ �{ �{ 
| | 2| P| `| t| �| �| �| �| �| �| �| �| }  } 2} D} T} f} v} �} �} �} �} �} �} �} 
~ ~ (~ 2~ >~ R~ b~ t~ �~ �~ �~ �~ �~ �~ �~  " < V d v � � � � � �     Jz         ����������P�`�p�����        q	�)K�"�3�        ���*                ��OR       �   [ C     ��OR          �[ �C ���������������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?�[�# ` p �p 0�0 � `�    \�# G	G	P( p( �( d\�# �* p) P( p( �( generic unknown error   �\�# �* �) P( p( �( iostream    iostream stream error    ]�# �* 0* ( p( �( system  3D-COAT preference.ini  Exchange    3D-CoatV3   Folder ..\MyDocuments\3D-CoatV3\Exchange not found! export.txt  File exists!    To import a new object? Start import!   d:\program files\maxon\cinema 4d r15\plugins\applink_cinema4dr15\source\applinkdialog.cpp   Start export!   open    3D-Coat.exe not found!  3D-Coat.exe is run! invalid string position string too long -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?���������������������������N���������������C}Ô%�I��}Ô%�I�TStop    obj output.obj  import.txt  
   [SkipImport]
   [SkipExport]
    write success! File    #Wavefront OBJ Export for 3D-Coat
  %d.%m.%Y  %H:%M:%S  #File created:  #Cinema4D Version:  Export object   Name    object. Material not found on   Default " has no UVW tag.
UV coordinates can't be exported. Object "    No selected objects!    [   ppp mv  ptex    uv  ref retopo  vox alpha   prim    curv    autopo  ]   d:\program files\maxon\cinema 4d r15\plugins\applink_cinema4dr15\source\applinkexporter.cpp  vertices
  # begin         v   # end    texture vertices
  vt  mtl mtllib  g    faces
 usemtl  f   /   newmtl  Ka 0.300000 0.300000 0.300000
  Kd  Ks  Ns 50.000000
   Tr 0.000000
    illum 2
    map_    d:\program files\maxon\cinema 4d r15\resource\_api\ge_dynamicarray.h          �?      ����������������������������N���������������C}Ô%�I��}Ô%�I�T����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?-DT�!	@-DT�!�?�`p#o.bad locale name �`�"G	G	�a#�'p$P909�9�9 :�99 9@bp#o.�bp#o.�]p!ios_base::badbit set    ios_base::failbit set   ios_base::eofbit set     ^p!$$�^� �#$    p^0"$$�D�D Q@T�S�T�U0LO�P ��?`� ,P4�BpF Q T�Q�T�U0K0NpP�Q�?P`� �#$    p    not found! Gathering of data...    vt  f       `_�"$$�D G QPT�S�T�U`L@O�P ��?�_� �#$    `   Wrong face in OBJ file! Nb Grp:     Nb faces:   .   Open file:  Parse file...   mtllib %s   g %s    v %lf %lf %lf   vt %lf %lf  vt %lf %lf %lf  Create objects...   V count:    Poly count:     Error on inserting phongTag. Object:    Selection   textures.txt     can not removed!   d:\program files\maxon\cinema 4d r15\plugins\applink_cinema4dr15\source\applinkimporter.cpp Open file   newmtl %s   Ns  Ns %lf  d   d %lf   illum   illum %d    Kd  Kd %lf %lf %lf  Ka  Ka %lf %lf %lf  Ks  Ks %lf %lf %lf  Ke  Ke %lf %lf %lf  map_Kd  map_Kd %s   map_Ks  map_Ks %s   displacement    displacement %f normalmap   Memory allocation error for material.   �b�"�'p$�8�8�8�8�8�9�8vector<T> too long  bad cast    �dy���=  �B    -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?���������������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?���������������������������N���������������C}Ô%�I��}Ô%�I�T�c�W�V`�p�����������d:\program files\maxon\cinema 4d r15\plugins\applink_cinema4dr15\source\applinkpreferences.cpp  icon_coat.tif   �cG	G	G	G	G	G	�a<dPc�c�e�e�d`dPa              �?                         -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�Td:\program files\maxon\cinema 4d r15\resource\_api\c4d_file.cpp -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?���������������������������N���������������C}Ô%�I��}Ô%�I�T�d`���������В �@�P�`�p��d�� �� �0�@�P�`�0e�� �� �0�@�P����d�� �� �0�@�P�`�|e�� �� �0�@�P����� �� �0�@�P�`������� �d:\program files\maxon\cinema 4d r15\resource\_api\c4d_gui.cpp  ~   Progress Thread 0%  %       -DT�!	@      Y@     �f@     @�@-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?���������������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�Td:\program files\maxon\cinema 4d r15\resource\_api\c4d_general.h       %s      -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�Td:\program files\maxon\cinema 4d r15\resource\_api\c4d_misc\memory\debugglobals.cpp %H:%M:%S     [%s %s L%d]    WARNING:    CRITICAL:   -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?���������������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?���������������������������N���������������C}Ô%�I��}Ô%�I�T�ep~0z    d:\program files\maxon\cinema 4d r15\resource\_api\c4d_baseobject.cpp   ����MbP?-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�Td:\program files\maxon\cinema 4d r15\resource\_api\c4d_resource.cpp #   M_EDITOR        -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�Tfp�-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�Td:\program files\maxon\cinema 4d r15\resource\_api\c4d_basebitmap.cpp   res     d:\program files\maxon\cinema 4d r15\resource\_api\c4d_misc\datastructures\basearray.h  -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?d:\program files\maxon\cinema 4d r15\resource\_api\c4d_pmain.cpp        -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?���������������������������N���������������C}Ô%�I��}Ô%�I�Td:\program files\maxon\cinema 4d r15\resource\_api\c4d_basetime.cpp        ����A  4&�kC �Ngm��C  4&�k�        ��������������       �       �-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T(f�� �G	G	    -DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?���������������������������N���������������C}Ô%�I��}Ô%�I�Td:\program files\maxon\cinema 4d r15\resource\_api\c4d_libs\lib_ngon.cpp        ���������������-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�T-DT�!	@-DT�!�?����������������������N���������������C}Ô%�I��}Ô%�I�Tw   pf��o.bad allocation  �f��o.g��o.Xg��o.       ���   ��   ��o   ���   ���   ��R   ���  ��  ��  �   ��7   ��d	  ���   �  $�p   8�P   ��   L�'   8�   ��   ��   h�   $�{   $�!   ���   ���   $��  ��   ��   ��   ��n   �a	  ���  ��   ��   L�   ��  ��   �    ��   ��   �   ��'  �@'  �A'  (�?'  @�5'  `�'  ��E'  ��M'  ��F'  ��7'  ��'  ��Q'  ��4'  �'  (�&'  4�H'  H�('  \�8'  p�O'  ��B'  ��D'  ��C'  ��G'  ��:'  ��I'  ��6'  ��='  �;'  $�9'  <�L'  P�3'  \�        f   t�d   ��e   ��q   ��   ��!   ��    �	   �h    �    ,�j   8�g   L�k   l�l   ��   ��m   ��   ��)   �   ��   ��   ��&   ��(   h�n   ��o   ��*           (�   $�   @    �   P s   ` t   p u   � v   � w   � 
   � y   � '   ��x   � z   � {   �    8�|         ��   L�   8   H�   X}   h~   x   ���   �i   ��p   �   ��   ��   ��   �   ���   �      ,$   D   ��"   d   x�   ��   ��   �   �   ��   �r   ��   �           permission denied   file exists no such device  filename too long   device or resource busy io error    directory not empty invalid argument    no space on device  no such file or directory   function not supported  no lock available   not enough memory   resource unavailable try again  cross device link   operation canceled  too many files open permission_denied   address_in_use  address_not_available   address_family_not_supported    connection_already_in_progress  bad_file_descriptor connection_aborted  connection_refused  connection_reset    destination_address_required    bad_address host_unreachable    operation_in_progress   interrupted invalid_argument    already_connected   too_many_files_open message_size    filename_too_long   network_down    network_reset   network_unreachable no_buffer_space no_protocol_option  not_connected   not_a_socket    operation_not_supported protocol_not_supported  wrong_protocol_type timed_out   operation_would_block   address family not supported    address in use  address not available   already connected   argument list too long  argument out of domain  bad address bad file descriptor bad message broken pipe connection aborted  connection already in progress  connection refused  connection reset    destination address required    executable format error file too large  host unreachable    identifier removed  illegal byte sequence   inappropriate io control operation  invalid seek    is a directory  message size    network down    network reset   network unreachable no buffer space no child process    no link no message available    no message  no protocol option  no stream resources no such device or address   no such process not a directory not a socket    not a stream    not connected   not supported   operation in progress   operation not permitted operation not supported operation would block   owner dead  protocol error  protocol not supported  read only file system   resource deadlock would occur   result out of range state not recoverable   stream timeout  text file busy  timed out   too many files open in system   too many links  too many symbolic link levels   value too large wrong protocol type �g��'p$*   C   ������������������������    r   a   rb  wb  ab  r+  w+  a+  r+b w+b a+b          
   !   "   2   *            #   3   +           -   0123456789abcdefghijklmnopqrstuvwxyz      !

					   0123456789abcdefghijklmnopqrstuvwxyz      A)!   0123456789abcdefABCDEF   	

   ��= �9 �3   ����?   ���9>   033�<   ����?   ���9>   033�<       ?  � ������?�              ?  � ������?�             �g��@h�-o.Unknown exception   Th�-o.csm�               �                      �?      �?3      3            �      0C       �       ��              fmod         D<�O��O�MMwM��O��?�h�@o.bad exception                                                                                                                                                                                                                                                                                     ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������k e r n e l 3 2 . d l l     FlsAlloc    FlsFree FlsGetValue FlsSetValue InitializeCriticalSectionEx CreateSemaphoreExW  SetThreadStackGuarantee CreateThreadpoolTimer   SetThreadpoolTimer  WaitForThreadpoolTimerCallbacks CloseThreadpoolTimer    CreateThreadpoolWait    SetThreadpoolWait   CloseThreadpoolWait FlushProcessWriteBuffers    FreeLibraryWhenCallbackReturns  GetCurrentProcessorNumber   GetLogicalProcessorInformation  CreateSymbolicLinkW SetDefaultDllDirectories    EnumSystemLocalesEx CompareStringEx GetDateFormatEx GetLocaleInfoEx GetTimeFormatEx GetUserDefaultLocaleName    IsValidLocaleName   LCMapStringEx   GetCurrentPackageId a m / p m   a / p      `   h   p   x   �   �   �   �	   �
   �   �   �   �   �   �   �   �   �   �                         (    0    8    @    H    P     X !   ` "   h #   p $   x %   � &   � '   � )   � *   � +   � ,   � -   � /   � 6   � 7   � 8   � 9   � >   � ?   � @   � A    !C   !D   !F   !G    !I   (!J   0!K   8!N   @!O   H!P   P!V   X!W   `!Z   h!e   p!   �  x!  �!  �!  �!  �!  �!  �!  �!	  �!  �!  �!  �!  "  "   "  ,"  8"  D"  P"  \"  h"  t"  �"  �"  �"  �"  �"  �"  �"   �"!  �""  �"#  �"$  #%  #&  #'  (#)  4#*  @#+  L#,  X#-  p#/  |#2  �#4  �#5  �#6  �#7  �#8  �#9  �#:  �#;  �#>  �#?   $@  $A  $C  $$D  <$E  H$F  T$G  `$I  l$J  x$K  �$L  �$N  �$O  �$P  �$R  �$V  �$W  �$Z  �$e  �$k  %l  %�  $%  0%  <%  H%	  T%
  `%  l%  x%  �%  �%  �%  �%  �%,  �%;  �%>  �%C  �%k  &  $&  0&  <&	  H&
  T&  `&  l&;  �&k  �&  �&  �&  �&	  �&
  �&  �&  �&;  �&  '  '  '	  ('
  4'  @'  L';  d'  t'	  �'
  �'  �'  �';  �'  �'	  �'
  �'  �';  (   (	   $(
   0(;   <($  L(	$  X(
$  d(;$  p((  �(	(  �(
(  �(,  �(	,  �(
,  �(0  �(	0  �(
0  �(4  �(	4  �(
4  )8  )
8  )<  ()
<  4)@  @)
@  L)
D  X)
H  d)
L  p)
P  |)|  �)|  �)�B   � ,   �)q   `    �)�   �)�   �)�   �)�   �)�   �)�   �)�    *�   *�   *�   $*�   0*�   <*C   H*�   T*�   `*�   � )   l*�   �*k   p !   �*c   h   �*D   �*}   �*�   p   �*E   �   �*G   �*�   �   �*H   �   +�   +�    +I   ,+�   8+�   p!A   D+�   �   T+J   �   `+�   l+�   x+�   �+�   �+�   �+�   �+�   �+�   �+�   �+�   �+K   �+�   �+�   �	   �+�   ,�   ,�    ,�   ,,�   8,�   D,�   P,�   \,�   h,�   t,�   �,�   �,�   �,�   �,�   �,�   �,�   �,�   �,�   � #   �,e   � *   �,l   � &   �,h   �
   -L   � .   -s   �   -�   (-�   4-�   @-M   L-�   X-�   X!>   d-�    !7   p-   �   |-N   � /   �-t   (    �-�   �-Z   �   �-O   � (   �-j   `    �-a   �   �-P   �   �-�   �-Q   �   �-R   � -    .r   � 1   .x   8!:   .�   �   `!?   $.�   4.S   � 2   @.y   � %   L.g   � $   X.f   d.�   � +   p.m   |.�   P!=   �.�   @!;   �.�   � 0   �.�   �.w   �.u   �.U   �   �.�   �.T   �.�        �.�   !6    /~       /V       /W   $/�   0/�   @/�   P/�       `/X        l/Y   H!<   x/�   �/�   �/v   �/�   0    �/[   x "   �/d   �/�   �/�   �/�   �/�    0�   0�   8     0\   �)�   ,0�   D0�   \0�   t0�   @    �0�   �0]    !3   �0z   h!@   �0�   (!8   �0�   0!9   �0�   H    �0^   �0n   P    �0_   !5   �0|   h     1b   X    1`   !4    1�   81{   � '   P1i   \1o   h1   x1�   �1�   �1�   �1�   �1�   �1F   �1p   a r     b g     c a     z h - C H S     c s     d a     d e     e l     e n     e s     f i     f r     h e     h u     i s     i t     j a     k o     n l     n o     p l     p t     r o     r u     h r     s k     s q     s v     t h     t r     u r     i d     u k     b e     s l     e t     l v     l t     f a     v i     h y     a z     e u     m k     a f     k a     f o     h i     m s     k k     k y     s w     u z     t t     p a     g u     t a     t e     k n     m r     s a     m n     g l     k o k   s y r   d i v   a r - S A   b g - B G   c a - E S   z h - T W   c s - C Z   d a - D K   d e - D E   e l - G R   e n - U S   f i - F I   f r - F R   h e - I L   h u - H U   i s - I S   i t - I T   j a - J P   k o - K R   n l - N L   n b - N O   p l - P L   p t - B R   r o - R O   r u - R U   h r - H R   s k - S K   s q - A L   s v - S E   t h - T H   t r - T R   u r - P K   i d - I D   u k - U A   b e - B Y   s l - S I   e t - E E   l v - L V   l t - L T   f a - I R   v i - V N   h y - A M   a z - A Z - L a t n     e u - E S   m k - M K   t n - Z A   x h - Z A   z u - Z A   a f - Z A   k a - G E   f o - F O   h i - I N   m t - M T   s e - N O   m s - M Y   k k - K Z   k y - K G   s w - K E   u z - U Z - L a t n     t t - R U   b n - I N   p a - I N   g u - I N   t a - I N   t e - I N   k n - I N   m l - I N   m r - I N   s a - I N   m n - M N   c y - G B   g l - E S   k o k - I N     s y r - S Y     d i v - M V     q u z - B O     n s - Z A   m i - N Z   a r - I Q   z h - C N   d e - C H   e n - G B   e s - M X   f r - B E   i t - C H   n l - B E   n n - N O   p t - P T   s r - S P - L a t n     s v - F I   a z - A Z - C y r l     s e - S E   m s - B N   u z - U Z - C y r l     q u z - E C     a r - E G   z h - H K   d e - A T   e n - A U   e s - E S   f r - C A   s r - S P - C y r l     s e - F I   q u z - P E     a r - L Y   z h - S G   d e - L U   e n - C A   e s - G T   f r - C H   h r - B A   s m j - N O     a r - D Z   z h - M O   d e - L I   e n - N Z   e s - C R   f r - L U   b s - B A - L a t n     s m j - S E     a r - M A   e n - I E   e s - P A   f r - M C   s r - B A - L a t n     s m a - N O     a r - T N   e n - Z A   e s - D O   s r - B A - C y r l     s m a - S E     a r - O M   e n - J M   e s - V E   s m s - F I     a r - Y E   e n - C B   e s - C O   s m n - F I     a r - S Y   e n - B Z   e s - P E   a r - J O   e n - T T   e s - A R   a r - L B   e n - Z W   e s - E C   a r - K W   e n - P H   e s - C L   a r - A E   e s - U Y   a r - B H   e s - P Y   a r - Q A   e s - B O   e s - S V   e s - H N   e s - N I   e s - P R   z h - C H T     s r     a f - z a   a r - a e   a r - b h   a r - d z   a r - e g   a r - i q   a r - j o   a r - k w   a r - l b   a r - l y   a r - m a   a r - o m   a r - q a   a r - s a   a r - s y   a r - t n   a r - y e   a z - a z - c y r l     a z - a z - l a t n     b e - b y   b g - b g   b n - i n   b s - b a - l a t n     c a - e s   c s - c z   c y - g b   d a - d k   d e - a t   d e - c h   d e - d e   d e - l i   d e - l u   d i v - m v     e l - g r   e n - a u   e n - b z   e n - c a   e n - c b   e n - g b   e n - i e   e n - j m   e n - n z   e n - p h   e n - t t   e n - u s   e n - z a   e n - z w   e s - a r   e s - b o   e s - c l   e s - c o   e s - c r   e s - d o   e s - e c   e s - e s   e s - g t   e s - h n   e s - m x   e s - n i   e s - p a   e s - p e   e s - p r   e s - p y   e s - s v   e s - u y   e s - v e   e t - e e   e u - e s   f a - i r   f i - f i   f o - f o   f r - b e   f r - c a   f r - c h   f r - f r   f r - l u   f r - m c   g l - e s   g u - i n   h e - i l   h i - i n   h r - b a   h r - h r   h u - h u   h y - a m   i d - i d   i s - i s   i t - c h   i t - i t   j a - j p   k a - g e   k k - k z   k n - i n   k o k - i n     k o - k r   k y - k g   l t - l t   l v - l v   m i - n z   m k - m k   m l - i n   m n - m n   m r - i n   m s - b n   m s - m y   m t - m t   n b - n o   n l - b e   n l - n l   n n - n o   n s - z a   p a - i n   p l - p l   p t - b r   p t - p t   q u z - b o     q u z - e c     q u z - p e     r o - r o   r u - r u   s a - i n   s e - f i   s e - n o   s e - s e   s k - s k   s l - s i   s m a - n o     s m a - s e     s m j - n o     s m j - s e     s m n - f i     s m s - f i     s q - a l   s r - b a - c y r l     s r - b a - l a t n     s r - s p - c y r l     s r - s p - l a t n     s v - f i   s v - s e   s w - k e   s y r - s y     t a - i n   t e - i n   t h - t h   t n - z a   t r - t r   t t - r u   u k - u a   u r - p k   u z - u z - c y r l     u z - u z - l a t n     v i - v n   x h - z a   z h - c h s     z h - c h t     z h - c n   z h - h k   z h - m o   z h - s g   z h - t w   z u - z a   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
         R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 4  
 -   i n c o n s i s t e n t   o n e x i t   b e g i n - e n d   v a r i a b l e s  
     D O M A I N   e r r o r  
     S I N G   e r r o r  
     T L O S S   e r r o r  
    
     r u n t i m e   e r r o r          ;   �1	   (2
   �2   �2    3   �3   �3    4   �4   �4   P5   �5   6   P6    7!   �7"   p9x   �9y   �9z   :�   0:�   8:R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
     R u n t i m e   E r r o r ! 
 
 P r o g r a m :     < p r o g r a m   n a m e   u n k n o w n >     . . .   
 
     M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y     m s c o r e e . d l l   CorExitProcess  ,"<%8"�!Sun Mon Tue Wed Thu Fri Sat Sunday  Monday  Tuesday Wednesday   Thursday    Friday  Saturday    Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec January February    March   April   June    July    August  September   October November    December    AM  PM  MM/dd/yy    dddd, MMMM dd, yyyy HH:mm:ss    S u n   M o n   T u e   W e d   T h u   F r i   S a t   S u n d a y     M o n d a y     T u e s d a y   W e d n e s d a y   T h u r s d a y     F r i d a y     S a t u r d a y     J a n   F e b   M a r   A p r   M a y   J u n   J u l   A u g   S e p   O c t   N o v   D e c   J a n u a r y   F e b r u a r y     M a r c h   A p r i l   J u n e     J u l y     A u g u s t     S e p t e m b e r   O c t o b e r   N o v e m b e r     D e c e m b e r     A M     P M     M M / d d / y y     d d d d ,   M M M M   d d ,   y y y y   H H : m m : s s          @    ީ@P�ީ(@P��P<@P��CT@P��Gl@P�3ML C _ A L L     L C _ C O L L A T E     L C _ C T Y P E     L C _ M O N E T A R Y   L C _ N U M E R I C     L C _ T I M E       	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ = ;     ;   =   C   _ . ,   _   .   �@�e+000         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          �      	         �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��log log10   exp pow asin    acos    exp10   atan    ceil    floor   modf    sin cos tan sqrt    (null)  ( n u l l )            EEE50 P    ( 8PX 700WP        `h````  xpxxxx          SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    TZ          �������             ��      �@      �               ���5�h!����?      �?  ccs UTF-8   UTF-16LE    UNICODE c c s   U T F - 8   U T F - 1 6 L E     U N I C O D E   sinh    cosh    tanh    atan2   fabs    ldexp   _cabs   _hypot  fmod    frexp   _y0 _y1 _yn _logb   _nextafter                    �?5�h!���>@�������             ��      �@      �        U S E R 3 2 . D L L     MessageBoxW GetActiveWindow GetLastActivePopup  GetUserObjectInformationW   GetProcessWindowStation \HE N U   pHE N U   �HE N U   �HE N A   �HN L B   �HE N C   �HZ H H   �HZ H I   IC H S   IZ H H   8IC H S   `IZ H I   �IC H T   �IN L B   �IE N U   �IE N A   JE N L   $JE N C   <JE N B   `JE N I   xJE N J   �JE N Z   �JE N S   �JE N T   KE N G   (KE N U   @KE N U   XKF R B   xKF R C   �KF R L   �KF R S   �KD E A   �KD E C    LD E L   DLD E S   `LE N I   |LI T S   �LN O R   �LN O R   �LN O N   �LP T B    ME S S   DME S B   dME S L   �ME S O   �ME S C   �ME S D   NE S F   $NE S E   LNE S G   pNE S H   �NE S M   �NE S N   �NE S I   �NE S A   OE S Z   <OE S R   XOE S U   �OE S Y   �OE S V   �OS V F   �OD E S   h E N G   �OE N U   �OE N U   a m e r i c a n     a m e r i c a n   e n g l i s h     a m e r i c a n - e n g l i s h     a u s t r a l i a n     b e l g i a n   c a n a d i a n     c h h   c h i   c h i n e s e   c h i n e s e - h o n g k o n g     c h i n e s e - s i m p l i f i e d     c h i n e s e - s i n g a p o r e   c h i n e s e - t r a d i t i o n a l   d u t c h - b e l g i a n   e n g l i s h - a m e r i c a n     e n g l i s h - a u s   e n g l i s h - b e l i z e     e n g l i s h - c a n   e n g l i s h - c a r i b b e a n   e n g l i s h - i r e   e n g l i s h - j a m a i c a   e n g l i s h - n z     e n g l i s h - s o u t h   a f r i c a     e n g l i s h - t r i n i d a d   y   t o b a g o   e n g l i s h - u k     e n g l i s h - u s     e n g l i s h - u s a   f r e n c h - b e l g i a n     f r e n c h - c a n a d i a n   f r e n c h - l u x e m b o u r g   f r e n c h - s w i s s     g e r m a n - a u s t r i a n   g e r m a n - l i c h t e n s t e i n   g e r m a n - l u x e m b o u r g   g e r m a n - s w i s s     i r i s h - e n g l i s h   i t a l i a n - s w i s s   n o r w e g i a n   n o r w e g i a n - b o k m a l     n o r w e g i a n - n y n o r s k   p o r t u g u e s e - b r a z i l i a n     s p a n i s h - a r g e n t i n a   s p a n i s h - b o l i v i a   s p a n i s h - c h i l e   s p a n i s h - c o l o m b i a     s p a n i s h - c o s t a   r i c a     s p a n i s h - d o m i n i c a n   r e p u b l i c     s p a n i s h - e c u a d o r   s p a n i s h - e l   s a l v a d o r   s p a n i s h - g u a t e m a l a   s p a n i s h - h o n d u r a s     s p a n i s h - m e x i c a n   s p a n i s h - m o d e r n     s p a n i s h - n i c a r a g u a   s p a n i s h - p a n a m a     s p a n i s h - p a r a g u a y     s p a n i s h - p e r u     s p a n i s h - p u e r t o   r i c o   s p a n i s h - u r u g u a y   s p a n i s h - v e n e z u e l a   s w e d i s h - f i n l a n d   s w i s s   u s     u s a   QU S A   $QG B R   4QC H N   @QC Z E   LQG B R   \QG B R   xQN L D   �QH K G   �QN Z L   �QN Z L   �QC H N   �QC H N   �QP R I   �QS V K   RZ A F   (RK O R   @RZ A F   \RK O R   tRT T O   h G B R   �RG B R   �RU S A   �OU S A   a m e r i c a   b r i t a i n   c h i n a   c z e c h   e n g l a n d   g r e a t   b r i t a i n   h o l l a n d   h o n g - k o n g   n e w - z e a l a n d   n z     p r   c h i n a     p r - c h i n a     p u e r t o - r i c o   s l o v a k     s o u t h   a f r i c a     s o u t h   k o r e a   s o u t h - a f r i c a     s o u t h - k o r e a   t r i n i d a d   &   t o b a g o   u n i t e d - k i n g d o m     u n i t e d - s t a t e s   A      A C P   O C P   6-�T�T�T�T�T�T�T�T�T�T�T U���Y�Y�Y�YZUUU U$U(U,U0U4U8UDU@HULU�PUTUXU����\U`UdUhUlUpU��tUxU|U�U�U�U�U�U�U�U�U�U�U�U�U�U�U�U�U�U�UV0VPVpV�V�V�V�VW4W\WxW�W�W�W�W�W�W�W�WX(XPXxX�X�X�XY0Y\Y�Y��__based(    __cdecl __pascal    __stdcall   __thiscall  __fastcall  __clrcall   __eabi  __ptr64 __restrict  __unaligned restrict(    new     delete =   >>  <<  !   ==  !=  []  operator    ->  ++  --  +   &   ->* <   <=  >   >=  ,   ()  ^   |   &&  ||  *=  +=  -=  /=  %=  >>= <<= &=  |=  ^=  `vftable'   `vbtable'   `vcall' `typeof'    `local static guard'    `string'    `vbase destructor'  `vector deleting destructor'    `default constructor closure'   `scalar deleting destructor'    `vector constructor iterator'   `vector destructor iterator'    `vector vbase constructor iterator' `virtual displacement map'  `eh vector constructor iterator'    `eh vector destructor iterator' `eh vector vbase constructor iterator'  `copy constructor closure'  `udt returning' `EH `RTTI   `local vftable' `local vftable constructor closure'  new[]   delete[]   `omni callsig'  `placement delete closure'  `placement delete[] closure'    `managed vector constructor iterator'   `managed vector destructor iterator'    `eh vector copy constructor iterator'   `eh vector vbase copy constructor iterator' `dynamic initializer for '  `dynamic atexit destructor for '    `vector copy constructor iterator'  `vector vbase copy constructor iterator'    `managed vector copy constructor iterator'  `local static thread guard'  Type Descriptor'    Base Class Descriptor at (  Base Class Array'   Class Hierarchy Descriptor'     Complete Object Locator'   CreateFile2 ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp       1#SNAN  1#IND   1#INF   1#QNAN  C O N O U T $       H                                                           H��h   RSDSe�p��h@���+�   D:\Program Files\MAXON\CINEMA 4D R15\plugins\applink_cinema4DR15\obj\Applink_Cinema4DR15_Win32_Release.pdb      4  4      L�        ����    @   �[           �[�[                d��[           �[ \�[    d�       ����    @   �[            ��0\           @\H\    ��        ����    @   0\            ��x\           �\�\H\    ��       ����    @   x\            А�\           �\�\�\H\    А       ����    @   �\            ��]           $]4]�\H\    ��       ����    @   ]��        ����    @   l]           |]P]                D��]           �]�]�]    D�       ����    @   �]`�       ����    @   �]           �]^    `�        ����    @   �]            |�4^           D^T^�]�]    |�       ����    @   4^            ���^           �^�^    ��        ����    @   �^          ��^           �^�^_(_D_    �       ����    @   �^|�              P   4^D�              @   �]`�              @   �]            0�t_           �_�_�^    0�       ����    @   t_    `      ���_           �_�_�^_(_D_    ��       ����    @   �_            ԓ`           (`4`�^    ԓ       ����    @   `    p      �d`           t`�`�^_(_D_    �       ����    @   d`            h��`           �`�`P]    h�       ����    @   �`            L�a           a a    L�        ����    @   al�       ����    @   Xa           ha<a a               �a�a<a a    ��       ����    @   ta           �a�a<a a    ��       ����    @   �a            ̔ b           b$b�a<a a    ̔       ����    @    b            ȑTb           dbtb�`P]    ȑ       ����    @   Tb            ���b           �b�btb�`P]    ��       ����    @   �b            ��b           cc�a<a a    �       ����    @   �b           HcTcpc    ��       ����    @   8c��        ����    @   �c           �cpc                ���c           �c�cTcpc    ��       ����    @   �c            ��d           d d    ��        ����    @   d            ��Pd           `dld d    ��       ����    @   Pd            h��d           �d�d�[    h�       ����    @   �d            L��[            ���d           ee    ��        ����    @   �d            ��De           Te`e�[    ��       ����    @   De            ���e           �e�e�d�[    ��       ����    @   �e            (��e           �e�e    (�        ����    @   �e            ���c             �<f           LfTf     �        ����    @   <f            ؝�f           �f�fP]    ؝       ����    @   �f            ���f           �f�fP]    ��       ����    @   �f            �g           ,g<g�fP]    �       ����    @   g            4�lg           |g�g�fP]    4�       ����    @   lg            X��g           �g�g<a a    X�       ����    @   �g            0�h           h$h    0�        ����    @   h            ��l]            (�hh           xh�hP]    (�       ����    @   hh             ��h           �h�hP]     �       ����    @   �h    �. /  � �' �z � � 0� P� p� �� �� �� �� � 0� P� p� �� �� �� �� � .�                             �,����    ����                  `i"�   pi   �i                            %+����    ����                  �i"�   �i   �i                            �>����    ����                  j"�    j   0j                            �J����    ����                  hj"�   xj   �j                            �/����    ����                  �j"�   �j   �j                            �I����    ����                  k"�   (k   8k                            �.����    ����                  pk"�   �k   �k                            �0����    ����                  �k"�   �k   �k                            �-����    ����                   l"�   0l   @l                            p
����    ����                  xl"�   �l   �l                            �����    ����                  �l"�   �l   �l                            �����    ����                  (m"�   8m   Hm                            �����    ����                  �m"�   �m   �m                            ����    ����                  �m"�   �m   �m                            �����    ����                  0n"�   @n   Pn                          �n   �n�n    h�    ����       �    ��    ����       �-          �n    oo�n�n    ��    ����       �    ȑ    ����       �    �-    Ho   To�n    (�    ����       -            |b����    ����                  po"�   �o   �o                            a����    ����                  �o"�   �o   �o                    ��    0p   <p�n    ؝    ����       *�    ��    ����       `�    ��    �p   �pXp�n    �    ����       E�    ��    �p   �pXp�n    4�    ����       {������"�   �p                       ����    ����    ����    �	    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    �         � ����    ����    ����    �!    ����    ����    ����    2#    ����    ����    ����    �#    ����    ����    ����    s&    ����    ����    ����    �'    ����    ����    ����    �)    ����    ����    ����    �3    ����    ����    ����15K5    ����    ����    ����    �?    ����    ����    ����    L    �K�K����    ����    ����     B    LAVA����    ����    ����I�I    ����    ����    ����A@J@@           �B����    ����                  Ls"�   \s   ls                   ����    ����    �����JK    �@    �s   �s�n     �    ����       l@    ����    ����    ����    mY    ����    ����    ����    /Z    ����    ����    ����    =[    ����    ����    ����    p�    ����    ����    ����    ˞    ����    ����    ����    v�    ����    ����    ����    ��    ����    ����    ����    D�����    P�����    ����    ����    ������    è����    ����    ����    ��        m�        |�    ����    ����    ����    թ    ����    ����    ����    ��    ����    ����    ����    '�    ����    ����    ����    ��    ����    ����    ����    ��    ����    |���    ����    ��    ����    ����    ����    ��    ����    ����    ����    h�    ����    ����    ����    ��    ����    ����    ��������    ����    ����    ��������    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    H    ����    ����    ����    }$    ����    ����    ����    n,    ����    ����    ����    �.    ����    ����    �����7�7    ����    ����    ����)B<B    ����    ����    ����    :n        lm����    ����    ����    �l    ����    ����    ����    Tr    ����    ����    ����    }�x         <z  � �y         \z P�                     �y �y 
z z ,z � � hz |z �z �z �z �z �z �z { { 2{ H{ Z{ j{ v{ �{ �{ �{ �{ �{ �{ 
| | 2| P| `| t| �| �| �| �| �| �| �| �| }  } 2} D} T} f} v} �} �} �} �} �} �} �} 
~ ~ (~ 2~ >~ R~ b~ t~ �~ �~ �~ �~ �~ �~ �~  " < V d v � � � � � �     Jz     � CloseHandle 
CreateToolhelp32Snapshot  'Process32First  )Process32Next �Module32First KERNEL32.dll  0ShellExecuteExA SHELL32.dll �IsDebuggerPresent qInterlockedIncrement  mInterlockedDecrement  @EnterCriticalSection  �LeaveCriticalSection  DeleteCriticalSection _Sleep <EncodePointer DecodePointer �WideCharToMultiByte �MultiByteToWideChar �GetStringTypeW  jGetLastError  QHeapFree  HRaiseException  �RtlUnwind �GetCommandLineA (GetCurrentThreadId  MHeapAlloc �GetSystemTimeAsFileTime fInitializeCriticalSectionAndSpinCount �GetCPInfo �UnhandledExceptionFilter  PSetUnhandledExceptionFilter SetLastError  #GetCurrentProcess oTerminateProcess  �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �GetStartupInfoW �GetModuleHandleW  �GetProcAddress  �IsProcessorFeaturePresent -GetDateFormatW  GetTimeFormatW  � CompareStringW  �LCMapStringW  nGetLocaleInfoW  �IsValidLocale GetUserDefaultLCID  aEnumSystemLocalesW  �GetStdHandle  �WriteFile }GetModuleFileNameW  mExitProcess �GetModuleHandleExW  , AreFileApisANSI VHeapSize  �IsValidCodePage �GetACP  �GetOEMCP  �FlushFileBuffers  �GetConsoleCP  GetConsoleMode  WGetFileType XReadFile  	SetFilePointerEx  #DeleteFileW �GetProcessHeap  |GetModuleFileNameA  <QueryPerformanceCounter $GetCurrentProcessId @GetEnvironmentStringsW  �FreeEnvironmentStringsW GetTimeZoneInformation  THeapReAlloc SetFilePointer  OutputDebugStringW  �LoadLibraryExW  �LoadLibraryW  /SetStdHandle  �WriteConsoleW VReadConsoleW  � CreateFileW �SetEndOfFile  �SetEnvironmentVariableA               ��OR    R�          H� L� P� �� j�   Applink_Cinema4DR15.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                              ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���P�d    .?AVGeDialog@@  d    .?AVApplinkDialog@@ d    .?AVerror_category@std@@    d    .?AV_Generic_error_category@std@@   d    .?AV_Iostream_error_category@std@@  d    .?AV_System_error_category@std@@    ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�Td    .?AVruntime_error@std@@ d    .?AVexception@std@@ d    .?AVfailure@ios_base@std@@  d    .?AVsystem_error@std@@  ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�Td    .?AVbad_cast@std@@  d    .?AVios_base@std@@  d    .?AV?$_Iosb@H@std@@ d    .?AV?$basic_ios@DU?$char_traits@D@std@@@std@@   d    .?AV?$basic_streambuf@DU?$char_traits@D@std@@@std@@ d    .?AV?$basic_istream@DU?$char_traits@D@std@@@std@@       d    .?AV?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    d    .?AV?$basic_istringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    d    .?AV?$basic_filebuf@DU?$char_traits@D@std@@@std@@   d    .?AV?$basic_ifstream@DU?$char_traits@D@std@@@std@@  d    .?AV_Facet_base@std@@   d    .?AVfacet@locale@std@@  d    .?AVcodecvt_base@std@@  d    .?AUctype_base@std@@    d    .?AV?$ctype@D@std@@ d    .?AV?$codecvt@DDH@std@@ ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�Td    .?AVCommandData@@   d    .?AVBaseData@@  d    .?AVApplinkPreferences@@    d    .?AVTriangulator@@  d    .?AVCTriangulator@TRIANGULATOR@@    ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�Td    .?AVSubDialog@@ d    .?AVGeUserArea@@    d    .?AVGeModalDialog@@ d    .?AViCustomGui@@        ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T      ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T       ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�Td    .?AVNeighbor@@  ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�Td    .?AVC4DThread@@ ���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�T���������������}Ô%�I��}Ô%�I�Td    .?AVbad_alloc@std@@ d    .?AVlogic_error@std@@   d    .?AVlength_error@std@@  d    .?AVout_of_range@std@@  ����d    .?AV_Locimp@locale@std@@       
       Copyright (c) 1992-2004 by P.J. Plauger, licensed by Dinkumware, Ltd. ALL RIGHTS RESERVED.                       �              �             �               3              �9               A                         �              �              �             �              �<              @>              2@      �<              @>              2@                     �              �             �        d    .?AVtype_info@@ N�@���Du�  s�   �     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       d    .?AVbad_exception@std@@ ��	����   8�.   4�L�L�L�L�L�L�L�L�L���P�P�P�P�P�P�P�.                                        	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 sqrt                            ��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                                                                                                                                                                                                                                                                                                   abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                                     abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                            ����            C       d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<==�<= =(=0=<=D=P=\=`=d=p=�=       �=�=�=�=�=�=�=�=�=�=�=> >0>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>d>�>�>�>??,?@?T?\?d?x?�?�!��                                   P�            P�            P�            P�            P�                          8�        ��X�                        �� �   �����	llllllllll    �����
                                                                  ?  �B�B    �p     ����    PST                                                             PDT                                                              �`�����        ����              �      ���������              �   LB   PB   @B   DB   D   D!   $D   TB   \B   lB   ,D   �B   �B   �B    �B   tB   |B   4D   �B   <D   DD   LD   TD   \D"   dD#   hD$   lD%   pD&   xD       �D        � 0                                                                                                                                                                                                                  �            �&  ����   :   Y   w   �   �   �   �     /  M  l  ����   ;   Z   x   �   �   �   �     0  N  m     ���5      @   �  �   ����             ����         �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                                                                                                                                                                                                                                                                                                                       �   080�021N1_1q1y1�1�1�1K2e2v2�2�2�2�2�2�2�2�23'3:3M3`3s3�3�3�3�3�3�3�344�4�4�455`5q5�5�5�516c6�6�67A7s7�7�7�7
8�8�8�8�8�8�9�9�9�9�9:!:A:U:g:x:�:�:�:�:�:�:";H;a;�;�;�;<8<J<[<o<�<h=y=�=�=�=�=>>P>b>t>�>�>�>�>�>�>??/?E?      8   z1V22D3X3�3�3�4�4�4�4�6�6�6�7,888`9�9 :E:�:�:�: 0    R1c1�1�1�1�12=2N2`2z2�2�2�2�2�263G3a3�3�3�3�3�304A4[4�4�4�4�4%5�5�5�56!6X6i6z6�6�6�6�6�677!7d7u7�7�7�7�7�7�7
88+8S8o8�8�8�8�8�899'9;9L9�9�9�9�9�9�9�9:B:S:e:m:~:�:�:�:�:�:;#;4;E;^;z;�;�;�;�;�;�;	<<.<B<V<g<x<�<�<�<=.=P=d=y=�=�=�=�=�=>>F>Z>~>�>Y?�?�?�?   @  �   r0�0�0�01!1)1C1T11�1�1�12t2�2�2�2�3�8�8�9�;�;*<g<{<�<�<�<�<�<==/=@=\=p=�=�=�=�=�=�=�=�=>">3>K>\>�>�>�>�>�>??0?A?h?�?�?   P  x  0?0d0{0�0�0�0�01:1P1b1j1{1�1�1�1�1�1�122.2G2X2m2�2�2�2�2�2�2�213B3T3\3m33�3�3�3�3�3�3 4"494N4w4�4�4�4�45*5?5S5d5|5�5�5�5�5�566(6<6X6l6�6�6�6�6�6�67-7E7Y7r7�7�7�7�7�7�7�788/8C8W8h8y8�8�8�8�8�8999=9Q9c9z9�9�9�9�9�9�9:#:8:I:Z:k:|:�:�:�:�:;%;-;>;P;\;w;�;�;�;�;�;�;<<*<><W<h<y<�<�<�<�<�<==(===E=Y=n=v=�=�=�=�=�=>'>8>`>w>�>�>�>�>??*?E?\?{?�?�?�?�?�?   `  l  0&0E0Y0t0�0�0�0�0�01 181L1h1}1�1�1�1�1�1�122.2B2V2j2~2�2�2�2�2�2�233*3?3G3[3s3�3�3�3�3�3	414H4]4�4�4�4�4�4�45.5M5a5|5�5�5�5�5�56+6F6]6|6�6�6�6�6�67'7F7^7r7�7�7�7�7�7�7�78&8:8N8b8{8�8�8�8�8�8�8�89#9+9?9W9z9�9�9�9�9�9:2:G:l:�:�:�:�:�:;;7;K;f;};�;�;�;�;<<0<G<f<z<�<�<�<�<�<=0=H=\=p=�=�=�=�=�=�=�=>$>8>L>e>�>�>�>�>�>�>�>�>??-?E?a?�?�?�?�?�? p  t  0020W0}0�0�0�0�0�0�01'1<1P1l1}1�1�1�1�1�12!252P2g2�2�2�2�2�2 33(3<3M3^3o3�3�3�3�3�3�3�34D4X4m4u4�4�4�4�4�4�4�45"565O5`5u5�5�5�5�5�5�5�56,6R6z6�6�6�6>7O7a7{7�7�7�7�7�7�7%898J8^8}8�8�8�8�8�899%979?9V9j99�9�9�9�9�9�9:":3:D:U:n:�:�:�:�:�:;;:;N;`;t;�;�;�;�;�;�;<<2<C<T<e<v<�<�<�<�<�<�<=#=j={=�=�=�=�=�=�=>>$><>P>l>}>�>�>�>�>�>�>
??4?S?q?�?�?�?�?�?�? �  4  
00&0B0c0~0�0�0�0�0�01-1?1G1[1t1�1�1�1�1�12 2U2f2x2�2�2�2�2�23 323:3N3c3k3�3�3�3�3�3�344-4B4V4o4�4�4�4�4�4�4�45.5B5z5�5�5�5�56#6W6h6z6�6�67-7>7P7X7i7{7�7�7�7�7�7�7�78&8?8T8e8v8�8�8�8�8�8�8�89*9C9p9�9�9�9�9�9::4:<:T:h:�:�:�:�:�:�:�:;#;4;F;N;c;t;�;�;f<�<�<�<2=L=`=p=�=�=�=6>S>�>?'?�?�?�? �  D  �0�0�0�011*1?1S1l1�1�1�1�1�1�1�1�122N2e2z2�2�2�2�2343K3`3t3�3�3�3�3�3�34#474O4f4�4�4�4�4�4�455.5?5X5i5z5�5�5�5�5�5�5 66"6;6�6�6�677$7,7=7R7f77�7�7�7�7�7�7	88+8<8H8l8�8�8�8�8�8�8�89989j9{9D:\:k:�:�:�:�:�:�:�:#;4;F;d;u;�;�;�;�;�;�;	<'<8<J<h<y<�<�<�<�<�<�<=4=E=W=p=�=�=�=�=�=�=�=�= >>>>>>>> >�?�? �  \   00D0U0}1�1�1�1>2�3�4�4�4�4�5@7�8�8�8�8�9�9�9�9�:0;�;�;�;�;�<:=�=5?Z?n?�?�?�?�?�?   �    0&0;0O0g0{0�0�0�0�0�081L1i1�1�1�1�1�162J2g2�2�2�23*323F3[3v3�3�3�3�3�344I4]4q4�4�4�4�4�4�45!585S5j5�5�5�5�5�56606D6�6�6�6�6�6�6�67f7z7�7�7�7P8�8�8�8-9U9z9�9�9�9�9�9:&:=:X:o:�:�:�:�:�:;!;5;I;p;�;�;�;�;�;�;<<3<G<b<y<�<�<�<�<�<�=�=�=>+>H>~>�>�>�>�>?2?a?}?�?�?�? �  �   0B0^0|0�0�0�0171�1�1252O2d2l2�2�2�2�23333S3h3p3�3�3�3�34 4445%5D5d5�5�5�6�6�6�6�7�7�7�7I8]8r8z8�8�8�8�8�8�8
9!9@9T9o9�9�9�9�9�9::C:u:�:�:�:�:F;~;�;&<�<�<==D=}=�=�=$>=>O>k>�>�>�>G?h?�?�?�?   �  �   0:0d0}0�0�0�0�0<1�1�1�12D2]2o2�2�2�23g3�3�3	4=4g4�4�4�4�4�4<5�5�5�56G6{6�6777K7S7g7{7�7�7�7�7�7�78+8F8]8�8�8�8�8�899 949I9Q9e9~9�9�9�9�9�9:,:W:k::�:�:�:�:;;6;�;<|<�<>>.>I>�>
?�?�?�?�?   �  h   0@0c0�0�0�0�0H3�326g6�6�67O7s7�9�:J;�;�;�;�;�;�;�;�;<)<G<^<}<�<�<�<�<==*=>=^=s=�=%>^>�>#?   �  �   �0O1c1x1�12o2�2�2�2�2�2�3�3�3�3�34 444H4c4z4�4�4�475[5�5�56:6W6�6�67'7;7�7�7�7<8\8u8�8�8�8�8�8�89 949H9c9z9�9�9�9�9�9
::0:G:\:p:�:�:�:�:�:; ;9;�>�>
??3?;?Q?h?�?�?�?�?�?   �   00Y0l0�0�0"161K1S1p1�1�1�1�1�1�1202D2X2l2�2313D3�3�3�45^5p5�5�5�5�56$6B6g6�8�8::*:�:�:�:�:�:�<�<�<�<�<q=>$>H>c>�?�?  �   &060�0�0V1f1�1�1�4�45555!5�5�5�5�5�56666!6�6�6�6�6�6�627]7�7�7�7�798_8�8�9:�:�:�:�:;;*;>;q;�;�;�;�;�<�<�<�<�<�<U=r=�=�=�=>a>u>�>�>?(?<?P?d?   \   181K1y1�1�12<2�2�2�23K3�3�4L6n6�67[8&:8:J;�;�;�;�;�;�;�;&<6<�<�<�<�=�=�>�>�?�?   0 d   1�1E2�2�4�435N5[5i5s5�5�5�5�5�566 6*6�667P7]7k7u7�7�7�7H<�<�<�<�<�<�<V=h=~>�>�>�>?&?4?A? @ \   Q0~0�0�0�0�0�0�1�1
22,212>2L2V2d2n2�2�8�8�9:�;�;8<@<�<�<�=�=�=>�>�>? ?g?m?�?�?   P 0   70�1�6	7+797J7\7g7�78�8�8J9�:�<�<�<=   ` �   �0�0�1�1�183B7H7N7T7d7�7�7�7[8|8�8�8�8�8$9d9�9�9�9:':Q:b:�:�:�:�:�:�:;;#;A;R;t;�;�;�;�; <<4<T<l<�<�<�<�<�<�< ===/=c=v=�=�=�=�=�=�=>$>D>d>�>�>�>�>�>$?6?D?V?t?�?�?�?�? p   0 0A0T0q0�0�0�0�01!111A1Q1d1�1�1�1�12$2D2d2�2�2�2�2353w3�3�3�344N4�4�4�4�45545d5�5�5�5�5�546R6m6�6�6�67$7D7d7�7�7�7�7848T8p8�8�8�8�89.9H9\9p9�9�9�9:D:h:�:�:�:;.;P;r;�;�;�;<<<`<�<�<�<!=4=d=�=�=�=�=>>!>1>A>Q>d>�>�>�>�>�>�>?$?Q?a?t?�?�?�?�?�?�?   �    0"020Q0d0�0�0�0�0141T1t1�1�1�1�12D2d2�2�2�2�2343T3t3�3�3�3�3444a4�4�4�4�45$5D5d5�5�5�5�56$6D6d6�6�6�6�67$7D7d7�7�7�7�7848T8q8�8�8�8�89919A9Q9a9t9�9�9�9�9�9:$:D:d:�:�:�:�:;6;N;x;�;�;�;�;<$<D<d<�<�<�<�<�<�<�<$=>=R=`=o=�=�=�=>>+>9>P>d>}>�>�>�>�>�>??4?T?t?�?�?�?�?   � �   0$0A0d0�0�0�0�01$1D1d1u1�1�1�1�1222Y2`2�2�2u3�3!494T4m4/5p5�5�5616Q6q6�6�6�6�6'7A7d7�7�7�7�7�78/8I8S8f8o8�8�8�8�89#9C9W9k9�9�9�9�9�9:":6:_:q:�:�:�:�:�:�:�:$;I;w;�;�;<O<�<�<='=Q=q=�=�=�=>7>g>�>�>�>?7?h?�?�?�?   � �   070d0�0�0�0101H1Y1�1'2Q2q2�2�2�2�2�2d3�3�3�4�45=5z5�5�5�56!6Q6�6�6�6717k7�7808J8b8z8�8�8�8�89W9y9�9�9�9�90:M:o:�:�:L;T;\;w;�;a<�<�<=h=�=�=�=�=>>>P>�>�>�>�>?P?�?�? � �   ;0{0�0�01u1�1�1�112e2�2�2�23K3�3�34�4'5V5^5f5�5�5!6�6�67,7N7b7t7�7�7�7+8m8�8�89f9�9�9�9:1:}:�:�:
;4;O;�;�;�;<*<L<`<�<�<�<�>�>�>�>J?   � �   =0]0v0�0�0�0 1a1�1�1�1!2Q2w2�2�2,343d3�34d4�45T5�5�5D6�6�647�7�7$8t8�89T9�9�9;:�:�:8;Y;�;<,<q<�<�<!=d=�=�=�=!>Q>�>�>-?m?�?�?�?   � �   0G0`0�0�0�0;1{1�1�1=2}2�2�2343a3�3�3414d4�4�455q5�5�5�56&6�6�67D7f7�7�7�7�7�7!8W88�8�8�89-9f9k9p9�9�9�9�9:w:�:�:9;�;3<�<�<�<�<�<�<�<�<�<�<�=>>>>> >$>(>,>�>�> ??8?A?d?�? � �   	00070?0m0�0�0�1�1�2�2c3�3�3444T4t4�4�4�4�4�45E5V5h5p5�5�5�5�5�5�5�56*6;6d6�6�6�6!7P7u7�7�7�7�7�718Q8l8�8�8�8�8!999Q9�9�9�9�9&:W:l:~:�:�:�:�:�:�:;;/;[;l;};�;�;�;<@<J<]<f<o<�<�<=D=y=�=>�>�>�>�>�>�>�>�>???A?_?{?�?�?   � �   /0D0t0�0�01d1|1�1�1�1�1�1�12202L2�2�2�23363g3�3454�4Y5{5'6:6�6�6+78$8l8s8�9:0:Q:t:�:�:�:;4;a;t;�;�;�;$<D<a<�<�<�<�<=G=q=�=�=�=�=$>D>d>�>�>�>�>?$?D?d?�?�?�?�?�?     |   010T0�0
1�12'2�2�23l3�3�3�4�4%5�5�5A6�6�6�67G7�7-8G8d8�8�89D9�9:7:T:p:�:;�;�;�;�;<|< ==�=>'>D>`>�>�>�?�?    �   0�0�0$1a1�1�1�1�1272d2�2�2�23E3a3t3�3�3�34!4D4a4�4�4�4�45!5G5w5�5�56!646T6t6�6�6�6�67!7@7E7J7O7d7�7�7�7�7�78D8^8�8�8�8�89T9�9�9:C:�:�:;T;t;�;�;<4<Q<d<�<�<�<=7=d=�=�=�=�=>G>t>�>�>�>!?1?D?d?�?�?�?�?�?     00$0D0d0�0�0�0�011"131H1\1t1�1�1�1�1�12"222T2n2�2�2�2�2�2343T3t3�3�3�3�3�34$4A4T4t4�4�4�4�4545`5�5�5�5�56 6A6Q6d6�6�6�647T7t7�7�7�7�78$8D8�8�8�8�89!959E9d9�9�9�9�9�9:G:�:�:�:;$;D;d;�;�;�;<$<A<T<z<�<�<�<�<�<�<3=s=�=�=>7>a>�>�>�>�>(?;?d?�?�?�?�?�? 0   080]0~0�0�0�01,1@1P1t1�1�1�12$2<2\2�2�2�2�233=3d3w3�3�3�3�3�3%4=4]4�4�4�4�4�45-5E5e5�5�5�5�56%6E6l66�6�6�6�6717D7d7�7�7�7�78$8D8d8�8�8�8�89$9D9a9q9�9�9�9:D:W:;3;�;�;�;�;�;;<\<p<�<�<�<�<�<=	==D=I=j=t=�=�=�=�=�=
>>2>j>�>�>�>+?3?8?B?G?Q?]?b?p?y?�?�?   @ �   0$0D0d0�0�0�0�0�0141T1q1�1�1�1$2I2l2�2�2�23343Q3d3�3�3�3�3�34!444Q4a4t4�4�4�4�4545^5�5�5�5�5�5616N6t6�6�6�6�67(7;7H9�9!:T:�:%;e;�;�;T<�<�<D=�=>8>k>>�>�>�>�>???f?�?�?�?�? P �   +0?0O0k0�0�0�0�0181h1|1�1�1�1242T2t2�2�2�23$3A3a3�3�3�3�34$4D4�4�4�4�4$5T5�5�5�5�56$6A6d6�6�6�6�6!7Z7�7�7�7$8A8g8�8�8�8�8A9`9x9�9�9�9:4:Q:t:�:�:�:	;&;T;k;�;�;�;�;<<O<j<�<�<�<�<=4=a=�=�=�=�=>Q>t>�>�>�>$?G?w?�?�?�? ` �   040T0t0�0�01:1e1y1�1�1�12!2A2a2�2�2�2333H3�3�3?4�4�4�4525d5�5�5�5�5!6q6�6�6�6747T7q7�7�7�78$8G8t8�8�8�8�8949g9�9�9�9:$:A:T:q:�:�:�:4;�;�;�;<4<o<�<�<=A=x=�=�=�=>/>I>g>�>}?�? p `   D0k0�0�2r5�56X6�6�8�8�8�8�8�89<9t9�9�9:::4:\:�:�:;$;G;�;�;;<t<�<�<�<'=a=�=�={>�>�? � �   �1�12$2D2a2�2�2�2�2343T3q3�3�3�344�45$5Q5t5�5�5�56!6D6T6�6�6�6�67$7Q7q7�7�7�7�7848T8�8�8�8�8919T9t9�9�9D:�:�:�:;4;T;t;�;�;�;<$<A<d<�<�<�<7=a=�=b>�>�>�>?u?�?�?�? � �   !0U0}0�0�0151u1�1�12%2e2�2�213b3�3�3�34Q4y4�4�4�4�45,5Q5y5�5�56W6�6�6�6-7m7�7�728b8�8�89R9�9�9:U:�:�:;E;u;�;�;5<�<�<�<%=V=�=�=%>e>�>�>%?u?�? � 0  0D0x0�0�0�0�01T1�1$2[2�2�2�2E3J3u3�3�3�3�3�3�3�3�34(4B4m4�4�4�4�4�4�455*5;5M5U5t5�5�5�5�5�5
6616E6e66�6�6�6�6�6�677+7=7E7d7x7�7�7�7�7�78!858U8o8�8�8�8�8�8�899+9U9d9p9�9�9�9�9�9�9�9:!:M:g:x:�:�:�:�:�:�:;";*;I;];};�;�;�;�;�;�;</<@<S<x<�<==>=�=�=�=�=�=><>P>p>�>�>�>�>�>U?f?w??�?�? � �   0050I0[0l0�0�0�0�011F1O1X1^1p1z1�1�1�1�122$2a2t2�2�2�2�23!343T3|3�3�3�3444r4�4�4�4545R5f5v5�5�5�56!616A6Q6a6t6�6�67'7T7q7�7�7�7�7878d8�8�8�8$979K9�9�9�9�9:1:T:t:�:�:�:;);Q;d;�;�;<<"<5<><Q<�<�<===1=s=�=�=>$>D>d>�>�>�>�>?$?A?T? � l   �0�0G1�1�1�122�2�3414D4a4t4�6�6�6�6�7�7�8�89"9h9�9�9:�:	<�<>=G=N=U=\=c=j=q=x=�=3>D>U>	?w?�?�?�? � �   !0G0�0�0�0�0�0�0�0�0�0�0�01*1B1R1y1�1�1W2�2�2�2�2�23=3E3�3�3�3�3�3�3�3�34,4?4F4Y4b4n4�4�4�4�4�4�4D5b5�5�5�5�5%6t6z6�6�6�6�6�6�67;7z7�7�7�7�7�7�7#898�8�8�8919Q9q9�9�9�9�9�9�<�<->e>U?�?�?   �     52`2�788888�:�:�:�= � p   �0�0�0%1e1�1�1%2b2�2�23B3u3�3�354r4�4�4525e5�5�5%6e6�6�6%7e7�78U8�8�8%9u9:�:>E>�>�>?:?U?p?�?�?�?�?     0040?0b0m0|0�0�0�0�0�0�0�01.141>1N1n1�34?4Q4a4�4
55"5*5?5\5q5}5�5�5676�6�6�6�6�6�67,787x7~78&8�8�8�8�8�8�8999.949:9A9I9O9�9�9�9�9�9�9�9g:l:u:�:�:#;K;Y;=#=<=C=K=P=T=X=�=�=�=�=�=�=�=�=�=�=�=2>8><>@>D>�>�>�>�>�>�>�>?/?a?h?l?p?t?x?|?�?�?�?�?�?�?�?  �   ]1�3�3�34A4�5o6�6�6�6�8�8�8�8�8�8�8�89'9E9L9P9T9X9\9`9d9h9�9�9�9�9�9*:5:P:W:\:`:d:�:�:�:�:�:�:�:�:�: ;;N;T;X;\;`;�<=c=�=�=�=�=�=�=�=�=�=�=�=�=�=>	>>>>>�>�?   �   060A0c0�0�0Y1`1�1�1B2�2�2�2�2|36�6y7�7r8�8�899�9�9�9�9�9�9:::*:5:=:J:T:z:�:�:�:�:;<;B;T;(=D=^=|=�=�=�=w>�>�>�?�?   0 �   03080�1�1�2�2�2383M3W3a3�3�3�3�3R4g4�4�45�5�5�5�5"6j6�67!7*727`8m8�8�8�8�;1<;<>J>r>�>�>�>�>�>�>�>�>�>#?V?e?l?�?�?�?�?�?�?�? @ <   |0�0�0�0�2�4�6�6�6T79�9b;�=�=8?C?c?n?�?�?�?�?�?�?   P 8  k0s0�0�0�0�193 44 4*4K4�4$56�6�6�6�6�6�6&7/7=7v77�7�7	9&989|9�9�:O;U;e;m;s;�;�;�;�;�;�;�;�;�;�;�;<<'<8<><D<K<T<Y<_<g<l<r<z<<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<=
====%=*=0=8===C=K=P=V=^=c=h=q=v=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>	>>>>!>'>/>4>:>B>G>M>U>Z>`>h>n>|>�>�>�>�>�>�>�?   `    $080h0�6�889u=   p    83   � �   @5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5q6�6]7v7�7�8�8999U9�9�9:::::?:E:K:V:\:�:�:�:�:�:�:�:;	;;.;4;O;Y;_;�;�<�<�<�<�<=>=Q=a=�=�=�=�=�=�=�=�=>%>1>8>A>Z>d>�>�>�>?x? � �   �0+1E1R1~1�1�1�1�1�1�1�1�1�12)222M2Y2_2j2x2~2�2�2�2�2�2�2�2�2�2�2�2�2.363I3T3Y3k3v3{3�3�3�3�3Y4p4}4�4�4�4�4�4�4�4�4 5#5(54595X5�5�5�5�516�6�6�6	7K7�7�8�8�8�8P9^9w9�9�9�9�9�9�9�9�9y:�:�;$<|<6=i=�=>^>p>�>?$?5?_?f?m?t?�?�?�?�?�?�?   � �   0Y0t0�1�1,292C2Q2Z2d2�2 33&393S3[3f3}3�3�3�3�3�3�3�3�3474q4�4�4T5�5�5�5(6�6�6�677`7z7�7�7�7�788+8P8l8�8�8�89*9C9T9�9�9�9�9�9o:�:;<�<==�=@?�?�?   � �   (030@0K0V0^0�0�011X1x1�1�1�182�2�2'373�4�6�6�7�7�7R8Y8l8�8�8�8�8�8�8�8�8�8�8�8�8�8�8999 9%9+959?9O9_9o9x9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::: :&:0:::M:R:(;I;N;   � d   s0�01�2�3N6T6Z6�6�6�6�6k7�7�7�7#8N8k8�8�8�8	9<9V9r9�9i:�:;";@;�;]<�<�<�<�<�=�=�=�>�>�?�?   � |   �0�0�0!1t1�1�1�2�263i3~3�3�3�34'4Z4u4�4�4�4�45L5^5�5�5�56*666�67�7�7�7'8�8�8>9 :C;J;�;�;�;<�<�<�<==�=i>�>�>   �    �5�5�>A?b?i?�?�?�?�? � �   22+272@2�2�2�2�23"3'3�4�4�4�4�4�4@5F5�6�67&7j7v7�7�7�7�7�7�7�788=8E8T8�8�8�8�8�8�8�8 99#9E9[9c9i9r9�9:T:]:l:x:�:�:�:�:�:�:;4;;;D;M;V;_;k;w;�;�;�;�;�;�;<<<<<<<<#<'<+</<;<Q<�<=�=�=�=�=f>{>�>     �    2�2a4g4�4�4�4�4S6}8�8�8�8�8�8�8�8�9�9�9�9�9�9:�;�;I<T<i<w<�<=="=/=7=?=G=O=X=a=i=u=}=�=�=�=�=�=�=�=�=�=�=H>N>�>�>�>3?9?@?F?^?t?�?�?�?�?�?�?    |    0000*020?0`0j0�0�0G2U2�2�2(343[3`3f3p3z3�3�3�3�3�3�3�5�5U6�6�677(74798�8H9�97;t;�;�;�<�<�<�<�<�=�=�=�>�>�>?     �   J0%1a1�1�1j2t3�3�3�3�344+404=4B4�46P6o6�6�6%717<8p8�8D9}9�9�9<:`:�:�;�;�;<'<�<�<�<==#=(=-=2=;=�=�=�=�=�=�=�=�=�=U>_>|>�>�> 0 �   �0!12!272M2U2]3�5�6�6|7�7�7�768H8Z8�8�:�;<<%<5<F<�=�=�=�=�=�= >>> >&>5><>L>R>X>`>f>l>t>z>�>�>�>�>�>�>�>�>�>�>�>�>�>@?X?q?   @ `   B0�0�1�1�1�1�1�1�2�2�2�2�2�233&383J3\3n3�3�3�3�6�67S7e7w7�7�7�7-9<9�9�9�9�9�9�=�=�=   P 0   �6�7�7A8_:;);�;�;�<�<1=>m>�>�>U?^?�?�? ` |   0\0�0Y1�1O2.3?3b3�3�3�3�384�4�4�4�4L5�5�5�5V6>8�8:<4<[<|<�<�<�<�<6=S=c=�=�=�=�=>T>d>}>�>�>�>?A?Q?c?�?�?�?�?�?   p �   
0�0�0?1N1m1~1�1�12�2�2�3�3�34424J4m4�4�4�4�4�4�45�5�5�5�5�5S6�6�6�6�677Z7p78�8�8�8�899'9�9�9�:1;=;�;�;�;<<�<=`=h=y=�=�=�>�>�?   � <   +30363=3�3@5T6b6|6�6�6�6�67�9:N:w:�:�:�:;}=�=�>�? � D   0)111�2k3w3444(4�4�4 5w5�6�6I8�8�8u9{9�9�9$:;:p:�:N>`>   � 4   �1�1�1�1�1�1�1�1�1�1�1�1�1�2�2�2�2W3�3�=�?�? � P   000&0=0h0}1�23�3�3�34f4�4�4�45[9l9�9�9�9�9�9�9D:X:�:;�;�;<�?�?   � p   0"0B0b0�0�0�0�01"1B1b1�1�1�1�12%2@2Q2a2q2�2�2�2�2�2�2�2�2�2�2�2�23333&3/383>3P3Z3h3}3�3�3�3�3�3   � h  \1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�233333 3$3L3P3T3X3\3`3d3094989L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 ::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;�=�=�=�=�=�=�=�=�=�=�=H?L?P?T?X?\?`?d?h?l?�?�?�?�?�?�?�?�? � �    00000000h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4�:�:�:p>t>   � \  `3d3h3l3p3�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666$6,646<6D6L6T6\6d6l6t6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7,747<7D7L7T7\7d7l7t7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888$848<8D8L8T8\8d8l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89999$9,949<9D9L9T9\9d9l9t9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9::::$:,:4:<:D:L:T:\:d:l:t:|:�:�:�:�:     h   034383<3P3T3X3\3`3d3h3l3p3t3x3|3�3�3`5d5h5l5p5t5�5�5�5 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6    �  $1,141<1D1L1T1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2,242<2D2L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444$4,444<4D4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�45555$5,545<5D5L5T5\5d5l5t5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666$6,646<6D6L6T6\6d6l6t6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7,747<7D7L7T7\7d7l7t7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888$8,848<8@8H8P8X8`8h8p8x8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 9999 9(90989@9H9P9X9`9h9p9x9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::: :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ==== =(=0=8=@=H=P=X=`=h=p=x=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>> >(>0>8>@>H>P>X>`>h>p>x>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???? ?(?0?8?@?H?P?X? 0 `   \:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;T<X<\<`<�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? @ �   $1(1P5\5h5t5�5�5�5�5�5�5�5�5�5�5�5666(646@6L6X6d6p6|6�6�6�6�6�6�6�6�6�6�6 777$707<7H7T7`7l7x7�7�7�7�7�7�7�7�7�7�7�788 8,888D8P8   P �   000$000<0H0T0`0l0x0�0�0�0�0�0�0�0�0�0�0�01 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�: ;�;�;�;�;�;�;�;�;�; <<(<,<<<@<H<`<p<t<�<�<�<�<�<�<�<�<�<�<�<�<�<== =$=(=,=4=L=P=h=x=|=�=�=�=�=�=�=�=�=�=�=�=>>,>0>@>D>H>L>T>l>|>�>�>�>�>�>�>�>�>�>�>�>�>�>??$?(?@?D?\?l?p?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   ` p   000$0(0,040L0\0`0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0 1111 181<1T1d1h1l1�1�1�1�1�1�1�1�1�1�1�1�1�1�122222$2<2L2P2`2d2h2l2t2�2�2�2�2�2�2�2�2�2�2�2�233333343D3H3L3T3l3p3�3�3�3�3�3�3�3�3�3�3�3 4444 484H4L4\4`4d4l4�4�4�4�4�4�4�4�4�4�4�4�4555,5<5@5P5T5X5`5x5�5�5�5�5�5�5�5�5�5�5�5�5�56 6$64686H6L6T6l6|6�6�6�6�6�6�6�6�6�6�6�6�6777(7,70747<7T7d7h7x7|7�7�7�7�7�7�7�7�7�7�7�7�78888$8<8L8P8`8d8t8x8|8�8�8�8�8�8�8�8�8�8l9�9�9�9�9�9�9�9:@:L:T:t:�:�:�:�:�:�:;$;H;T;\;|;�;�;�;�;�;<<,<P<\<d<�<�<�<�<�< ===4=X=d=l=�=�=�=�=�=>>><>`>l>t>�>�>�>�>�>�>�>�>�>�>�>�>�>�>?? ?4?<?D?L?P?X?l?|?�?�?�?�?�?   p �   00$0,04080@0T0\0p0x0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�001P1p1�1�1�1�1�1282X2x2�2�2�2�2�2�2 333$3(3D3H3X3|3�3�3�3�3�3�3�3�3�3�3484X4x4�4�4�4�45 5,5H5T5`5�5�5�5�5 6 6@6`6�6�6�6�6�6�6 7 7@7`7�7�7�7�7�7�7�78(8H8   � d   @0D0H0L0d0�0�0�0�0h1�1�1�1(2D2`2|2�2�203�3�34L4l4�4�4�4�4�5�5�5�5�5h7�7�7�7(: =�=�=>4>X>   � \  00X0`0 4 4$40484<4@4D4H4L4P4T4X4\4h4l4p4t4x4|4�4�4 6X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<==$=D=P=T=X=\=x=|=�=�=�=�=�=�=�=�=�=�=�=>>�>�>�>�>�>????$?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    