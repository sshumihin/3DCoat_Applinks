MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       `�r$�x!$�x!$�x!���!%�x!-��!�x!-��!��x!u!!�x!$�y!D�x!-��!s�x!-��!%�x!-��!%�x!Rich$�x!                        PE  L %LM        � !	  \  �      .�     p                         �                              �� Q   �� <                            0 T6  �q                            `� @            p \                          .text   �[     \                   `.rdata  r   p  t   `             @  @.data   �:   �     �             @  �.reloc  �A   0  B   �             @  B                                                                                                                                                                                                                                                                                                                                                                                        U���V��H�Q`V�ҡ��U�H�E�IdRj�PV�у���^]� ���������̡��P�BlQ��Y�U��j�hCId�    PQV�p�3�P�E�d�    ��u��BR �N�E�    ��q��A �N$�E��A� �ƋM�d�    Y^��]����������������U��j�hqId�    PQV�p�3�P�E�d�    ��u���q�N$�E�   蒪 �N�E� �B ���E�������Q �M�d�    Y^��]���������U���T  �p�3ŉE�Wj j�@ ����u_�M�3��^� ��]�V������PWǅ����(  �d@ ����   ������Qj�T@ �����   ������RPǅ����$  �(@ ���}   ������P������h  Q�"� ������h  R蕾 ���������P�I �@��u�+�$    ��/t��t������H��\uꍴ����V�j� hrV�"� ����u.������PW�? ���8���W� p^3�_�M�3��]� ��]ËM�^3͸   _�H� ��]���������j j j�r �����U��j�h�Id�    P��`SVW�p�3�P�E�d�    ��E�P�M�Q3ۋ��E�   �]��Z 9]��&  �M���� ���B�P`�M�Q�]��҃��E�Pj�M܍~Q���E��E P�M��E��� �U�R�M��E��� �M��E��Q� ���H�Al�U�R�E��Ћ��Q�Jl�E�P�]��у�hDr�M�臧 �U�R�M��E��ש �M��]���� �E�SP袶 �����L  ���Q�J`�E�P�ы��B�PdSj��M�h4rQ�ҍE�P�E��� ���Q�Jl�E�P�]��у�S����Q ���B�P`�M�Q�ҡ��H�AdSj��U�hrR�ЍM�jQ�E��� �����B�Pl�M�Q�E�]��҃� S8]�t~hr�M������E�P�E��%� ���Q�Jl�E�P�]����� SSh8h�   �E��� ���E��E�;�t	���b�  �3��U�WR�Ȉ]���  h�  ���#Q �S�E�P���E�   �]���� �M��E�����茦 �M�d�    Y_^[��]� ��������U���SVW��j�~W�E�3�P�E�   �]��*� jW�M�Q���E�   �]��� jW�U�R���E�   �]��Z jW�E�P���E�   �]��Y jW�M�Q���E�   �]��Y jW�U�R���E�   �]��rY j
W�E�P���E�
   �]��Y j	W�M�Q���E�	   �]��BY jW�U�R���E�   �]��*Y j�E�   �]�W�E�P���Y jW�M�Q���E�   �]��:� jW�U�R���E�   �]���X _^[��]������������U��j�h�Jd�    P���   SVW�p�3�P�E�d�    ����t ����   h�r�M��Y� ��l���3�P�]��� �M�QP�U�R�E��� ���~$P���E�褦 �M��E�訤 ��l����]�蚤 �M��E�����苤 �^@�#� �E�SW�E�   �"� ������  �E�P���,� P�M��E��� Sj�M�Q�M��E��� ���M��E��E��*� ���B�Pl�M�Q�E��҃�8]�t'�E�P�E�����謵 ��3��M�d�    Y_^[��]�Sh�r�M��G����M�Q�~j���E��#D ���B�Pl�M�Q�E��҃�h�r�M��� h�r��l����E���� ��4���j	P�E�致 ��l���QP��P���R�E�	�� �M�QP�U�R�E�
�m� �� ��P����E��;� ��4����E��,� ��l����E��� �M��E��� �E�jP趱 ���M���tQ�M��ã Pj���E��EC �M��OShPr�E���P�E���� ���H�Al�U�R�E��Ѓ�Sh�r�M������M�Qj���E���B �M܋��B�PlQ�E��҃�Sj����A jj���A jj���A jj���A Sj
���A jj	���kA jj���`A Sj���VA Sh�r�M������E�Pj���E��gB ���Q�Jl�E�P�E��у�Sj���A �M�W�۹ �M��� �M��E��ǡ �U�R�N$苢 P�M��E��N� �M�Sj�E�P�E��{� ���M��E��E�艡 ���Q�Jl�E�P�E��у�8]�t'�U�R�E������� ��3��M�d�    Y_^[��]ËM�j�~W�Ƶ �M��>� ���E�   �]�H�A`�U�R�Ѓ��M�Qj�U�R���E��= SSP�E�P���E��iP ���Q�Jl�E�P�E��ы��B�Pl�M�Q�E��ҡ��E�   �]�H�A`�U�R�Ѓ��M�Qj�U�R���E��*= SSP�E�P���E���O ���Q�Jl�E��E�P�ы��B�Pl�M�Q�E��҃�h���h   �Sjh���h   �Sj���E�   �]��^: P�E�P���bL SSj���E�   �]���9 P�M�Q���Q� SSj���E�   �]���9 P�U�R���0� SSj���E�   �]��9 P�E�P���� h���h   �Sjh���h   �Sj
���E�
   �]���9 P�M�Q����K �E�	   �]�SSj	���S9 P�U�R��跊 SSj���E�   �]��29 P�E�P��薊 SSj���E�   �]��9 P�M�Q���u� ���E�   �]�B�P`�M�Q�҃��E�Pj�M�Q���E��; SSP�U�R���E��ON ���H�Al�U�R�E��Ћ��Q�Jl�E�P�E��у�SS�E�   �]�j���|8 P�U�R����� h�  ����H �E�P�E������� ���   �M�d�    Y_^[��]�����������U��j�h�Jd�    P��0VW�p�3�P�E�d�    ���@ ��   訯 �E��E�P�O$�E�    � P�M��E�腝 j j�M�Q�M��E�豯 �Mċ��E��Ý ���B�Pl�M�Q�E� �҃���t���/����M���W蓵 �M�蛯 �E�P�E������+� ���M�d�    Y_^��]��������U��j�h�Kd�    P��   SVW�p�3�P�E�d�    ��3ۉ]��F@   �����E����   ����   ����  ���H�A`�U�R�Ћ��Q�JdSj��E�hrP�эU�R�E�   ��� ���H�Al�U�R�E��������� SSh8h�   ���i� ��,�E�E�   ;�t	����  �3���VW���E������:�  �`  �MQ�U�R���E�   �]��<N 9]�>  h�  ���F �-  �=� SSh8j$���� ��;�t�@   ��X�X�X�X�3���VW���E�������F  ���H�A`�U�R�Ѓ��M�Qj�Uؿ   R�Ή}��]8 ���H�Al�U�R�E��Ѓ�Sj���5 ��t7Sh�r�M���������Q�R S�E�P�M�Q�E��}��҃��E��u�]�E��E�   t���H�Al�U�R�Ѓ�8]�  �����S����   ���Q�JP�E�P�ы����B��H  S�SV�ы�S���B�PTV�M�WQ��j<��L���SP襰 ��0��L���QǅL���<   ��P�����T���ǅX����r��\�����d���ǅh���   ��l����Tq��ueSh�r�M�������U�R�E��z� ���H�Al�U�R�E����0h�r�M������M�Q�E��I� ���B�Pl�M�Q�E��҃����H�Al�U�R�E������Ѓ��   �M�d�    Y_^[��]� ������������V��V臫 ���    ^�������������U��V��������Et	V�پ ����^]� �������������������������������U����UV��H�ApVR�Ѓ���^]� ��������������U���V��H�Q`V�ҡ��H�U�ApVR�Ѓ���^]� �����   �Q��Y���������������U������P�M�P��P�P�P�P �P�P�P,�P(�X$���Q�P�I�H�M��P�Q�P�I�H�M��P�Q�P�I�H �M��P$�Q�P(�I�H,]� ���U��M�U�A�
�E��A�J���A$�J����A�
�A�A�J���A(�J���X�A�
�A�A �J���A,�J���X�A�J�A�J���B�I$���X�A�J�A�J���B�I(���X�A �J�A�J���A,�J���X�A�J�A�J���B �I$���X�A�J�A�J���B �I(���X�A �J�A�J���A,�J ���X �B$�I�A�J(���B,�I$���X$�A�J(�A�J$���B,�I(���X(�A �J(�A�J$���A,�J,���X,]���U��U��t�M��t�E��tPRQ�@� ��]������������U��j�h�Kd�    P��SVW�p�3�P�E�d�    3ۉ]�]��E�M�Q�M�]��E؉]܉]�� �}S�U�R�E�P���E��^ �M���]��A� ;�t}�����   �JX�E�P�ы���;�t_�����   �PT���ҋ����   �M�RQPV�ҋ�����   ��U�R�E������Ѓ��ƋM�d�    Y_^[��]� �����   �
�E�P�E������у�3��M�d�    Y_^[��]� ������������U��j�hLd�    P�� SVW�p�3�P�E�d�    3ۉ]��]�]�E�M�Q�   �M��}��Eԉ]؉]��] �MS�U�R�E�P�E��( �M����E��
� ;�t\�����   �JH�E�P�ы��u���B�H`V�ы��B�HpVW�ы����   ��M�Q�E�   �]��҃��C���H�u�Q`V�ҡ��H�QdSj�h�rV�ҡ����   ��U�R�}��]��Ѓ��ƋM�d�    Y_^[��]� �U��j�h/Ld�    P��SV�p�3�P�E�d�    3ۉ]�]��E�M�Q�M�]��E؉]܉]��6 �MS�U�R�E�P�E�� �M���]���� ;�tJ�����   �J8�E�P�ы������   ��M�Q�E������҃��ƋM�d�    Y^[��]� �����   ��U�R�E������Ѓ�3��M�d�    Y^[��]� ����U��j�hkLd�    P�� SV�p�3�P�E�d�    3��u��u�u�E�M�Q�M��u��Eԉu؉u��C �MV�U�R�E�   P�]��]��
 ��t�����   �J�E�P�у���u2ۍM��u���� ��tK�����   �P<�M�Q���]�����   ��U�R�E��������E���M�d�    Y^[��]� �����   �
�E�P�E��������E���M�d�    Y^[��]� �������U��j�h�Ld�    P��SV�p�3�P�E�d�    3ۉ]�]��E�M�Q�M�]��E؉]܉]��& �MS�U�R�E�P�E��� �M���]���� �����   �E�P;�t7�J@�ы�u�H��P���N���   ��V�U�R�E������Ѓ����u�
�V�V�E�������у��ƋM�d�    Y^[��]� ���������U��j�h�Ld�    P�� SV�p�3�P�E�d�    3ۉ]��]�]�E�M�Q�M��E�   �Eԉ]؉]��/ �MS�U�R�E�P�E��� �M����E���� ;�tC�����   �JL�E�P�ыu��P���� �����   ��M�Q�E�   �]����(�uS���Z� �����   ��U�R�E�   �]��Ћƃ��M�d�    Y^[��]� �����U��j�h�Ld�    PQSVW�p�3�P�E�d�    ���H�AP�Uj3�R�}��Ћ��Q����H  WFWV�Ћ�j�E��Q�JTVP�EP��N��$;�~�]��$    �U��P��衚 G;�|�M�Q蓰 ���B�Pl�MQ�E������҃��M�d�    Y_^[��]� ���U��j�h Md�    P��SVW�p�3�P�E�d�    ���H�A`�U�R�Ћ��Q�Jd3�Wj��E�h�rP�ы��B�PP�M�jQ�}��ҋ���H��H  WFWV�ҋ�j�E��Q�JTVP�E�P��N��8;�~�]�U��P��諙 G;�|�M�Q蝯 ���B�Pl�M�Q�E������҃��M�d�    Y_^[��]� �������������U��Q�ESVW���   3�3�3�3ۃ��M�|#�@|�O���A�	�d$ p����u�E�M�;�}�@|��_�^�[��]� �����U��j�h�Md�    P��   SV�p�3�P�E�d�    3ۉ]���H�u�Q`V�]��ҡ��H�QdSj�h8sV�҃��E�]��E�   ��
�j  �$�p0 Sh4s�M��i����E�P���E�   �b  ���Q�Jl�E�P�]����&  Sh0s�M��/����U�R���E�   �mb  �U���  Sh(s�M������M�Q���E�   �Eb  ���B�Pl�M�Q�]�����  Sh$s��p����������p���P���E�   �b  ���Q�Jl��p���P�]����  Sh s�M������U�R���E�   ��a  �U��H  Shs��P����_�����P���Q���E�   �a  ���B�Pl��P���Q�]����  Shs�M������E�P���E�   �]a  ���Q�Jl�E�P�]�����   Shs�M�������U�R���E�   �#a  �U��   Shs�M������M�Q���E�	   ��`  ���B�Pl�M�Q�]����}Sh�r��`���������`���P���E�
   �`  ���Q�Jl��`���P�]����=Sh�r��@����C�����@���R���E�   �~`  ��@������H�AlR�]��Ѓ����Q�J`�E�P�ы��B�PdSj��M�h�rQ�ҡ��H�QV�E�   �ҋ��Q�R0�M�QPV�ҡ��H�Al�U�R�]��Ѓ�(�ƋM�d�    Y^[��]� �I �- �- �- %. h. �. �. / 5/ l/ �/ ����U��j�h9Nd�    PQSVW�p�3�P�E�d�    ���}�3��   �G�7�w�w�w�w�_�u��C�3�s�s�s�s�G@�w0�w4�wD�w<�w8�GX�wH�wL�w\�wT�wP�Gp�w`�wd�wt�wl�wh���   �wx�w|���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   �E�97t	W�l� ���7�w�w�w�w93t	S�Q� ���G0�3�s�s�s�s90t	P�3� ���GH�w0�w4�wD�w<�w890t	P�� ���G`�wH�wL�w\�wT�wP90t	P��� ���Gx�w`�wd�wt�wl�wh90t	P�֩ �����   �wx�w|���   ���   ���   90t	P諩 �����   ���   ���   ���   ���   ���   90t	P�z� �����   ���   ���   ���   ���   ���   �ǋM�d�    Y_^[��]����������������U��j�h�Nd�    PQSVW�p�3�P�E�d�    ��u��E�   �� ���   3��E�9t	W�� ����_�_�_�_���   �E�9t	W辨 ����_�_�_�_�~x�E�9t	W蜨 ����_�_�_�_�~`�E�9t	W�z� ����_�_�_�_�~H�E�9t	W�X� ����_�_�_�_�~0�E�9t	W�6� ����_�_�_�_�~�]�9t	W�� ����_�_�_�_�E�����9t	V�� ����^�^�^�^�M�d�    Y_^[��]�U��j�h�Od�    P��(  SVW�p�3�P�E�d�    ���}���H�A`�U�R�Ћ��Q�Jdj j��E�hXsP�ы��B�P`��|���Q�E�    �ҡ��H�Adj j���|���hLsR�ЋMQ�����R�E��G P��|���P��<���Q�E��/\  �U�RP�E�P�E��\  ��H���Q�Jl��<���P�E��ы��B�Pl�����Q�E��ҡ��H�Al��|���R�E��Ћ��Q�Jl�E�P�E��ы]���B�H`��S����e�V�ы��B�Pp�M�VQ�҃����/����u�~ �E�    �e  3����H�A`�U�R�Ћ��Q�Jdj j��E�h�rP�ы��B�P`�M�Q�E�	�ҡ��H�Adj j��U�hHsR�Ћ��Q�J`��\���P�E�
�ы��B�Pdj j���\���hHsQ�ҡ��H�A`�U�R�E��Ћ��Q�Jd��@j j��E�hDsP�у��F�D8j0j jj �Q�U��$�E�R�  ���؋F�D8j0j j�j Q��L����$P�E���� ���E�F�8j0j j�j Q��l����$Q�E���� P�U�R��,���P�E��Z  ��\���QP������R�E���Y  �MQP������R�E���Y  �M�QP�����R�E���Y  ��HSP������P�E��Y  �M�QP������R�E��Y  ���Q�Rp�M�QP�E��ҡ��H�Al������R�E��Ћ��Q�Jl������P�E��ы��B�Pl�����Q�E��ҡ��H�Al������R�E��Ћ��Q�Jl������P�E��ы��B�Pl��,���Q�E��ҡ��H�Al��l���R�E��Ћ��Q�Jl��L���P�E��ы��B�Pl�M���@Q�E��ҡ��H�Al�U�R�E����E�
���Q�Jl��\���P�ы��B�Pl�M�Q�E�	�ҡ��H�Al�U�R�E��ЋM���B��Q�H`���܉eS�ы��B�Pp�M�SQ�ҋM��������E�@��;F�E�������}�]���H�A`�U�R�Ћ��Q�Jdj j��E�hXsP�ы��B�P`�M�Q�E��ҡ��H�Adj j��U�h<sR�ЋMQ��l���R�E��� P�E�P��L���Q�E��W  �U�RP�E�P�E��oW  ��H���Q�Rp�M�QP�E��ҡ��H�Al�U�R�E��Ћ��Q�Jl��L���P�E��ы��E��B�Pl��l���Q�ҡ��H�Al�U�R�E��Ћ��Q�Jl�E�P�E��ы��B�H`��S����eV�ы��B�Pp�M�VQ�҃����[���S���#������H�Al�U�R�E������Ѓ��M�d�    Y_^[��]� ����U��j�h\Rd�    P��  SVW�p�3�P�E�d�    ���}���H�A`������R�Ћ��Q�Jdj j�������htsP�ы��B�P`�����Q�E�    �ҡ��H�Adj j������hLsR�Ћu�F,P������Q�E��� P�����R��(���P�E��U  ������QP�U�R�E��U  ��H���H�Al��(���R�E��Ћ��Q�Jl������P�E��ы��B�Pl������E�Q�ҡ��H�Al������R�E��ЋM���B��Q�H`���܉eS�ы��B�Pp�M�SQ�҃�������3�9]�]�  ���H�A`������R�Ћ��Q�Jdj j�������h�rP�ы��B�P`��x���Q�E�	�ҡ��H�Adj j���x���hHsR�Ћ��Q�J`������P�E�
�ы��B�Pdj j�������hHsQ�ҡ��H�A`������R�E��Ћ��Q�Jd��@j j�������hpsP�у��Fj0�<[j �j��D8�j �E�Q��(����$R�|� ���E��F�D8���j0j ��jj Q�]썅����E��E��$P�G� ���E�F�8j0j j�j Q�������$Q�E��� P������R��x���P�E��eS  ������QP��H���R�E��MS  �M�QP��H���R�E��8S  ��x���QP��h���R�E�� S  ��H�M�QP��X���R�E��S  ������QP��x���R�E���R  ���Q�Rp�M�QP�E��ҡ��H�Al��x���R�E��Ћ��Q�Jl��X���P�E��ы��B�Pl��h���Q�E��ҡ��H�Al��H���R�E��Ћ��Q�Jl��H���P�E��ы��B�Pl��x���Q�E��ҡ��H�Al������R�E��Ћ��Q�Jl�����P�E��ы��B�Pl��@��(���Q�E��ҡ��H�Al������R�E��Ћ��Q�Jl������P�E�
�ы��B�Pl��x���Q�E�	�ҡ��H�Al������R�E��ЋM����Q�J�Q`���ĉe�P�E��ҡ��H�U��IpR�E�P�ыM���������B�P`������Q�ҡ��H�Adj j�������h�rR�Ћ��Q�J`�E�P�E��ы��Bj j�hHs�M�Q�Pd�ҡ��H�A`������R�E��Ћ��Q�Jdj j�������hHsP�ы��B�P`��X���Q�E��ҡ��H�Ad��@j j���X���hpsR�Ѓ��N�Dj0j j�Dj Q��h����$R�E���� ���E�F�D�D��j0j ��jj Q�]��������E��E��$Q��� ���E��Vj0j �E��|j�j Q�������$P�� P��X���Q������R�E���O  ������QP������R�E���O  �M�QP�����R�E��O  �M�QP������R�E��O  ��H�M�QP������R�E� �O  ������QP������R�E�!�mO  ���Q�Rp�M�QP�E�"�ҡ��H�Al������R�E�!�Ћ��Q�Jl������P�E� �ы��E��B�Pl������Q�ҡ��H�Al�����R�E��Ћ��Q�Jl������P�E��ы��B�Pl������Q�E��ҡ��H�Al������R�E��Ћ��Q�Jl������P�E��ы��B�Pl��h�����@Q�E��ҡ��H�Al��X���R�E��Ћ��Q�Jl������P�E��ы��B�Pl�M�Q�E��ҡ��H�Al������R�E��ЋM��Q���e����B�H`��W�ы��B�Pp�M�WQ�ҋM���������H�A`��h���R�Ћ��Q�Jdj j���h���h�rP�ы��B�P`�M�Q�E�#�ҡ��H�Adj j��U�hHsR�Ћ��Q�J`�E�P�E�$�ы��B�Pdj j��M�hHsQ�ҡ��H�A`�����R�E�%�Ћ��Q��@j j�hps�����P�Jd�у��Fj0j �|[�j��D8�j Q��x����$R�E�&�~� ���E�F�D8���j0j ��jj Q�]��������E��E�'�$P�I� ���E��F�8j0j j�j Q�������$Q�E�(�� P�����R������P�E�)�gL  �M�QP������R�E�*�RL  �M�QP�����R�E�+�=L  �M�QP��8���R�E�,�(L  ��H�M�QP��X���R�E�-�L  ��h���QP��h���R�E�.��K  ���Q�Rp�M�QP�E�/�ҡ��H�Al��h���R�E�.�Ћ��Q�Jl��X���P�E�-�ы��B�Pl��8���Q�E�,�ҡ��H�Al�����R�E�+�Ћ��Q�Jl������P�E�*�ы��B�Pl������Q�E�)�ҡ��H�Al�������E�(R�Ћ��Q�Jl������P�E�'�ы��B�Pl��x�����@Q�E�&�ҡ��H�Al�����R�E�%�Ћ��Q�Jl�E�P�E�$�ы��B�Pl�M�Q�E�#�ҡ��H�Al��h���R�E��ЋM���B��Q�H`�����e�W�ы��B�Pp�M�WQ�ҋM�������N|�E�<��u  ���B�P`�M�Q�ҡ��H�Adj j��U�h�rR�Ћ��Q�J`�E�P�E�0�ы��B�Pdj j��M�hHsQ�ҡ��H�A`��(���R�E�1�Ћ��Q�Jdj j���(���hHsP�ы��B�P`��H���Q�E�2�ҡ��H�Ad��@j j���H���hpsR�Ѓ��Fj0�|[	j �j��D8�j �E�3Q��8����$Q��� ���E�F�D8���j0j ��jj Q�]��������E��E�4�$R��� ���E��F�8j0j j�j Q�������$P�E�5�� P��H���Q������R�E�6��H  ��(���QP������R�E�7��H  �M�QP������R�E�8�H  �M�QP�����R�E�9�H  ��H�M�QP��8���R�E�:�H  �M�QP��X���R�E�;�vH  ���Q�Rp�M�QP�E�<�ҡ��H�Al��X���R�E�;�Ћ��Q�Jl��8���P�E�:�ы��B�Pl�����Q�E�9�ҡ��H�Al������R�E�8�Ћ��Q�Jl������P�E�7�ы��B�Pl������Q�E�6�ҡ��H�Al������R�E�5�Ћ��Q�Jl������P�E�4�ы��B�Pl��@��8���Q�E�3�ҡ��H�Al��H���R�E�2�Ћ��Q�Jl��(���P�E�1�ы��B�Pl�M�Q�E�0�ҡ��H�Al�U�R�E��ЋM���B��Q�H`�����e�W�ы��B�Pp�M�WQ�ҋM�������E�N|�@;E�E������}���B�P`�M�Q�ҡ��H�Adj j��U�htsR�Ћ��Q�J`�E�P�E�=�ы��B�Pdj j��M�h<sQ�ҋv,������VP�E�>�\� P�M�Q������R�E�?�GF  �M�QP��8����@R�]��1F  ��H���Q�Rp�M�QP�E�A�ҡ��H�Al��8���R�]��Ћ��Q�Jl������P�E�?���E�>���B�Pl������Q�ҡ��H�Al�U�R�E�=�Ћ��Q�Jl�E�P�E��ы]���B�H`��S����eV�ы��B�Pp�M�VQ�҃�������S����������H�Al�U�R�E������Ѓ��M�d�    Y_^[��]� �U��j�h�Sd�    P���   SVW�p�3�P�E�d�    ����HH�U���  j h�  R�Ћ}��j j�ωE��$	 j j�ωE��	 ���Q�J`���E�P�}��у��E�    ���4  �~ �*  ��\����8n ��0���R�E��� ��聟 P��\����E��p ��0����E��n ���H�A`�U�R�Ћ��Q�Jdj j��E�h�sP�у��U�R��\����E���o ���H�Al�U�R�E��Ћ��Q�J`�E�P�ы��B�Pdj j��M�h�rQ�ҡ��H�A`�U�R�E��Ћ��Q�Jdj j��E�h�sP�у�,�E���0���R��\����Ո �M�Q���E��n P�U�R�E�P�E��dC  �M�QP�U��R�]��QC  ���Q�Rp�M�QP�E�	�ҡ��H�Al�U�R�]��Ћ��Q�Jl�E�P�E��ы��B�Pl�M�Q�E��҃�,��0����E��Hm ���H�Al�U�R�E��Ћ��Q�Jl�E�P�E��ы]��S���e�����B�H`W�ы��B�Pp�M�WQ�҃����2���S���������\����E� ��l ��]���H�A`�U�R�Ћ��Q�Jdj j��E�h�rP�ы��B�P`�M�Q�E�
�ҡ��H�Adj j��U�h�sR�Ѓ�(�����   �M�Bx�E���P�M�Q�U�R��A  �M�QP�U�R�E���A  ���Q�Rp�M�QP�E��ҡ��H�Al�U�R�E��Ћ��Q�Jl�E�P�E��ы��B�E�
�MċPlQ�ҡ��H�Al�U�R�E� �Ћ��Q�B`��0S�����eW�Ћ��Q�Jp�E�WP�у��������S�������U�}RWS���"����}� t�E��MPQWS���������B�P`�M�Q�ҡ��H�Adj j��U�h�sR�Ћ��Q�J`�E�P�E��ы��B�Pdj j��M�hLsQ�ҋEP�M�Q�E��� P�U�R�E�P�E��{@  �M�QP�U�R�E��i@  ��H���Q�Rp�M�QP�E��ҡ��H�Al�U�R�E��Ћ��Q�Jl�E�P�E��ы��E��B�Pl�M�Q�ҡ��H�Al�U�R�E��Ћ��Q�Jl�E�P�E� �ы��J�Q`��S���ĉeP�E�ҡ��H�U�IpR�E�P�у����V������B�P`��L���Q�E    �ҡ��H�Adj j���L���h�rR�Ћ��Q�J`��x���P�E��ы��B�Pdj j���x���h�rQ�҃�(�} �E��E    �  �}� ��  �~ ��  ���   �M�������   ����� ���   �ȋBx�Ћ��Q�Rp��x���QP�ҡ��H�I j ��L���R��x���P�у����_  ���B�P`�M�Q�ҡ��H�Adj j��U�h�rR�Ћ��Q�J`�E�P�E��ы��B�Pdj j��M�h�sQ�ҍ�x���P�M�Q�� ���R�E��'>  �M�QP�� ���R�E��>  ��@���Q�Rp�M�QP�E��ҡ��H�Al�� ���R�E��Ћ��Q�Jl�� ���P�E��ы��B�Pl�M�Q�E����E����H�Al�U�R�Ћ��Q��S���ĉe�EP�B`�Ћ��Q�E�RpP�M�Q�҃����������H�Ip��L���R��x���P�у����B�P`�����Q�ҡ��H�Adj j������h�sR�Ћ��Q�Rp�E�P�����Q�E��ҡ��H�Al�����R�E��ЋO|�U�� �<� �E    ��  �]�����    ���H�A`�U�R�Ћ��Q�Jdj j��E�hHsP�ы��B�P�M�Q�E��ҋ��Q�M�Q�J0P�E�P�ы��B�Pl�M�Q�E��ҋG4�N�ÍDP��<���Q�%� �E���B�P�M�Q�E��ҋ��Q�MQ�J0P�E�P�ы��B�Pl��<�����@Q�E��҃��}� ��   �\ ��   ���H�A`�U�R�Ћ��Q�Jdj j��E�h�sP�ы��B�P�M�Q�E��ҋ��Q�M�Q�J0P�E�P�ы��B�Pl�M�Q�E��ҋGL�N�ÍDP��h���Q�7� �E���B�P�M�Q�E��ҋ��Q�MQ�J0P�E�P�ы��B�Pl��h�����@Q�E��҃��E�O|�U@��;��E�����]���H�A`�U�R�Ћ��Q�Jdj j��E�h�rP�ы��B�P�M�Q�E��ҋ��Q�M�Q�J0P�E�P�ы��B�Pl�M�Q�E��ҋ��Q��(S���ĉe�EP�B`�Ћ��Q�E�RpP�M�Q�҃���������E�O|��U@;E�E��������H�A`�U�R�Ћ��Q�Jdj j��E�h�sP�ы��B�P`�M�Q�E��ҡ��H�Adj j��U�h<sR�ЋMQ�� ���R�E� �� P�E�P��<���Q�E�!�9  �U�RP��h���P�E�"�l9  ��H���Q�Rp�M�QP�E�#�ҡ��H�Al��h���R�E�"�Ћ��Q�Jl��<���P�E�!�ы��E� �B�Pl�� ���Q�ҡ��H�Al�U�R�E��Ћ��Q�Jl�E�P�E��ы��B�H`��S�����eW�ы��B�Pp�M�WQ�҃����U���S���������H�Al��x���R�E��Ћ��Q�Jl��L���P�E� �ы��B�Pl�M�Q�E������҃��M�d�    Y_^[��]� ������������U��j�h�Td�    P��  SVW�p�3�P�E�d�    ����H�A`��`���R�E�    �Ћ��Q�Jdj j���`���hHsP�э�`���R�EP�M�Q�E��7  ���B�Pl��`���Q�E��ҋE�]��$PS�M�Q���C������B�P`�M�Q�ҡ��H�Adj j��U�h�rR�Ћ��Q�J`�E�P�E��ы��B�Pdj j��M�hHsQ�ҡ��H�E���p����A`R�Ћ��Q�Jdj j���p���hHsP�у�<�E�j0j jj Q�U��$R�E��q� �����E�j0j jj Q�E��$P�E��P� ���E�E�j0j jj Q��P����$Q�E��+� ��p���RP��4���P�E�	�s6  �MQP�����R�E�
�^6  �M�QP������R�E��I6  W�E�P������P�76  ��H�M�QP�����R�E��6  �����H�A�U�R�E��Ћ��Q�J0WP�E�P�ы��B�Pl�����Q�E��ҡ��H�Al������R�E��Ћ��Q�Jl������P�E��ы��B�Pl�����Q�E�
�ҡ��H�Al��4���R�E�	�Ћ��Q�Jl��P���P�E��ы��B�Pl�M�Q�E��ҡ��H�E��Al�U�R�Ћ��Q�Jl��p���P�E��ы��B�Pl�Mă�@Q�E��ҡ��H�Al�U�R�E��ЋM���B��Q�H`�����eW�ы��B�Pp�M�WQ�҃����c����Eh�  PS����������~  h�  P��(���Q���6�����D����E��'^ ��M��]��^ ���M�U�R�E��(� ��D���QW��(���RP�E�诬 ���M��E��^ �M��]��^ ���H�A`�U�R�Ћ��Q�Jdj j��E�hHsP�ы��B�P`�M�Q�E��ҡ��H�Adj j��U�h�sR�ЍMQ�U�R�E�P�E��3  �E��M�QP�U�R�3  ��@���Q�Rp�M�QP�E��ҡ��H�Al�U�R�E��Ћ��Q�Jl�E�P�E��ы��B�Pl�M�Q�E��ҡ��H�Al�U�R�]��Ћ��Q�J`�E�P�ы��B�Pdj j��M�h�rQ�҃�,�E�P��D����E�� ^ �M�QP�U�R�E���2  �����H�U��E�R�A�Ћ��Q�J0WP�E�P�ы��B�Pl�M�Q�E��ҡ��H�Al�U�R�E��Ћ��Q�Jl�E�P�]��ыU���H��(R�Q`�����eW�ҡ��H�Ap�U�WR�Ѓ����������D����E��\ ��(����E��|\ ���Q�Jl�E�P�E� �ы��B�Pl�MQ�E������҃��M�d�    Y_^[��]�$ ������U��j�h}Ud�    P���   SVW�p�3�P�E�d�    ��M��K[ ���H�A`�U�R�E�    �Ѓ��M�Q�M�   S�U�R�E��f�  P��D����]��W[ ��D���P�M��E��T] ��D����]��[ ���Q�Jl�E�P�E��ы��B�Pl�M�Q�E� �ҋM����D���P�� P�M��E��] ��D����E� �<[ ���Q�J`�E�P�ы��B�Pdj j��M�h�sQ�҃��E��E�P�M��l\ ���Q�Jl�E�P�E� �у��U�R�M��[ P�E��ݦ ���H�Al�U�R�E� �Ѓ��p^ �E�h1D4ChCD4C�E����x� Pj S�M�Q���^ ��u;�U�R�E��I^ ���M��E�    �E������`Z 3��M�d�    Y_^[��]� �~ �E    ��  �F�M���<��B�P`�M�Q�ҡ��H�A`��p���R�E��Ћ��Q�Jdj j���p���h�rP�ы��B�P`�M�Q�E�	�ҡ��H�Adj j��U�htR�Ѓ�,�����   �Bx���E�
��P�M�Q��P���R�-/  ��p���QP��4���R�E��/  ���Q�Rp�M�QP�E��ҡ��H�Al��4���R�E��Ћ��Q�Jl��P���P�E�
�ы��B�Pl�M�Q�E�	�ҡ��H�Al��p���R�E��ЋM����B��0Q�H`���܉e�S�ы��B�Pp�M�SQ�҃����������H�A`�U�R�Ћ��Q�Jdj j��E�h�sP�ы��B�@p�M�Q�U�R�E��Ћ��Q�Jl�E�P�E��ыU���� R���e�܋H�Q`S�ҡ��H�Ap�U�SR�Ѓ�������h�  W���r�����tL���Q�B`���܉e�S�Ћ��Q�Bdj j�h�sS�ЋM��U��h4  h@  WQR���B���h�  W��������tJ���H�Q`���܉e�S�ҡ��H�Qdj j�h�sS�ҋE��M��h�	  hD  WPQ����������B�P`��`���Q�ҡ��H�Adj j���`���h�sR�Ћ��Q�Rp�E�P��`���Q�E��ҡ��H�Al��`���R�E��ЋM����B�� Q�H`�����e�W�ы��B�Pp�M�WQ�҃����%������H�A`�U�R�Ћ��Q�Jdj j��E�h�sP�ы��B�@p�M�Q�U�R�E��Ћ��Q�E��Jl�E�P�ыU���H�� R�Q`�����e�W�ҡ��H�Ap�U�WR�Ѓ����������Q�J`�E�P�ы��B�Pdj j��M�h�sQ�ҡ��H�Ip�U�R�E�P�E��ы��B�Pl�M�Q�E��ҋE����Q�� P�B`�����e�W�Ћ��Q�Jp�E�WP�у���������U�R���������H�Al�U�R�E��ЋE@��;F�E�=����M��Y �M�Q�E� �1Y ���M��E�    �E������HU �   �M�d�    Y_^[��]� ���������������U��j�h�Wd�    P��  SVW�p�3�P�E�d�    �ى�����hG  �c� �K ���� ��������  �������T ���H�A`�U�R�E�    �Ѓ��u�M�Qj�U�R���E��/�  P��(����E��T ��(���P�������E��V ��(����E��ZT ���Q�Jl�E�P�E��ы��B�Pl�M�Q�E� �ҋ}����(���P���ʄ P�������E���U ��(����E� ��S ���Q�J`��`���P�ы��B�Pdj j���`���h<uQ�҃��E���`���P�������U ���Q�Jl��`���P�E� �у���������R ���B�P`�M�Q�E��҃��E�Pj�M�Q���E����  P��(����E���R ��(���R�������E�	��T ��(����E��%S ���H�Al�U�R�E��Ћ��Q�Jl�E�P�E��у�h0u��(����WR ��(���R�������E�
�T ��(����E���R �������R ���H�U��E�R�A`�Ѓ��M�Qj�U�R���E��*�  P��(����E��R ��(���P�������E��T ��(����E��UR ���Q�Jl�E�P�E��ы��B�Pl�M�Q�E��҃�h$u��(����Q ��(���P�������E���S ��(����E���Q �M�Q�������R P�E��� ���B�Pl�M�Q�E��҃��E�P�������R P�E�趝 ���Q�E��E؋JlP�у��U�R�������NR P�E�脝 ���H�Al�U�R�E������Ũ��UЍM�� uQ�]ԍ����R��H���ٕ���P�荍d���ٕ ���QٝH�����x���ٕ$���ٕL���ٕP���ٕd���ٕh���ٝl������������   ���   �щE�j P���E���} �����   �M苐�   �҅���  �fT �E�h1D4ChCD4C�E����n� Pj j������P���{T ��uz�M�Q�E��:T ��3��u싂�   ���   �M�Q�E��҃��u荍�����E��4P �������E� �%P �������E������P 3��M�d�    Y_^[��]� j h�r�M��^����E�P�M�Q�������E��P ���ԉečM�QPR�E��`%  �����������B�Pl�M�Q�E��ҡ��H�Al�U�R�E��Ѓ�j h�r�M������M�Q�U�R�������E��2P ���̉ečU�RPQ�E���$  ����葾�����H�Al�U�R�E��Ћ��Q�Jl�E�P�E��у�j h�r�M��t����U�Rj j���E��1�  P�E�P���e������̉ečU�RPQ�E��n$  �����������H�Al�U�R�E��Ћ��Q�Jl�E�P�E��у�j j�����  P�U�R�������P�E�腚 ���H�Al�U�R�E��ЋM���R j hu�M�趢��j hu�M��E�裢��������E�Q��������N P�U�R��`���P�E��#  �M�QP�����R�E��#  P�E� ��� ���H�Al�����R�E��Ћ��Q�Jl��`���P�E��ы��B�Pl�����Q�E��ҡ��H�Al�U�R�E��Ћ��Q�Jl�E�P�E��у�0�,Q �E�h1D4ChCD4C�E�!���4� Pj j������R���AQ ��u6�E�P�E�� Q �M�3�Q�u��E���P ���M�u��E���  ��������B�P`��D���Q�҃�3�Wh�t�M��E�"�K������H�Ip��D���R�E�P�E�#�ы��B�Pl�M�Q�E�"�ҋE���P����D����̉e�R�>������׻���   ��4�����0�����,���Pǅ,����  ��@�����<�����8����N ��Wh�r�M�譠��Wh�t�M��E�$蛠����,���Q�����h�tR�E�%�/ P�E�P��`���Q�E�&�!  �E�'�U�RP�����P�!  ��$P��D����E�(�R������Q�Jl�����P�E�'�ы��B�Pl��`���Q�E�&�ҡ��H�Al�����R�E�%�Ћ��Q�Jl�E�P�E�$�ы��B�Pl�M�Q�E�"�ҋE���P����D����̉e�R������芺��Wh�r�M�蜟��Wh�t�M��E�)芟����� P�����Q�E�*�� P�U��E�+R��`���P�   �M�QP�����R�E�,�x   �� P��D����E�-�E������H�Al�����R�E�,�Ћ��Q�Jl��`���P�E�+�ы��B�Pl�����Q�E�*�ҡ��H�Al�U�R�E�)�Ћ��Q�Jl�E�P�E�"�ыU���R����D����̉e�P�������~����M�Q���C���Wj���	�  �M�{�{�����������   ���   ��\����҅��{  蓖 �����   ��\����M苒�   P�ҋ������   �B�ω}���=�  �	  ���Q�J`�����P�ы��B�Pdj j������h�tQ�҃������   �Bx���E�.��P�����Q������R��  P�E�/�� ���H�Al������R�E�.�Ћ��Q�Jl�����P�E�"�у��������������B�P`�����Q�E�0�ҡ��H�Adj j������h�tR�Ѓ������   �Bx���E�1��P�����Q������R�7  P�E�2蝔 ���H�Al������R�E�1�Ћ��Q�Jl�����P�E�0�у������� ��  ���BH���   h�  ��V�у�P��p����  j�������w  j ��p����J  ���E�    �,� ���u�����  �����   �P����=�  ��  hF  h�  V��诰�����{  j ���E�   �G� ������  h�  V�E�P��謱�����Q�J�E�P�E�7�у�����   W��������  �M��� ������   ���$    �d$ �����   �P����=)  ��   �����   �Bx���ЍM�Q���  ��tu���� ��X���R������Q3�V�ȉE���� ��tO�	��$    ��������F;�X������������t���J��@;�X���~�M���X���R������PV�� ��u������   �B(���Ћ����/�����������9j ��p����  ���B�Pl�M�Q�E�0�ҋu��������   �B(���Ћ��E����.����������9 ��   ���B�P`�M�Q�ҡ��H�Adj j��U�h�tR�Ѓ������   �� �����@|�U�R�E�8�Ћ��Q�Jl�E�P�E�0�ы���JT�Q,j P�҃�����
  ������Q���,� �荕d���ٕd���Rٕh���h�  ٝl����������E�9�m�  ���������������E�0��  �}� ��   ������ �E�    ��   ��    3�9{~a���$    �S����� ���   �ȋBx�Ћ������Uȋ�������   �Bx�Ћ��Qj VP�B �Ѓ���t1G;{|��s�������Uȋ<���|jjjV���  ��t�C�<��E�@;������E��Z������QH�u����  j h�  V�Ћ��QHj ��������  h�  V�Ћ��QH�E����   h�  V�Ћ��QH�E����   h�  V�Ћ���h�����(�}�;�t(}+�PW��T����  �jj��+�QP��T�����  3���~-�u�����I �3�;V��X�����@����;ǉL��|�u��}�������P��蝴����l���������;�t(}+�PW�������,  �jj��+�QP�������  ��H���R���'� P��x���P��p���Q裪���E��E����E�3Ƀ��E��E��)  �u����������G����F��    �U�م|����������H�T8��؅p����E��H������H����]̋]��E��H�؅t������H������H����]��E��H�؅x������H������H��]ЉY���]ԋ]�م|����Y�H��������L؅p����E��H���������]̋U��E��H�؅t������H���������]��E��H�؅x������H��������UЉQ���]ԋU�م|����Q�H؅p����E��H������ȍW������H���]̋U��E��H؅t������H�����H���]��E��H؅x������H�����H��UЉQ���]ԋU�م|����Q�H�������W�؅p�����E��H�����H��ٝT����E��H؅t������H�����H���]��E��H؅x������H�����H���]�مT����]̋U��E���]ЋU��E��Q�]ԋUԃ�0���Q������Mċ�����;M���   ������I������D�+�U�+�م|����������H��ȃ���؅p����E��H������H���ٝT����E��H�؅t������H������H����]��E��H�؅x������H������H����]�مT����]̋}��E��9�]Ћ}��E��y�]ԋ}ԉy�f�����l����܋� �����������;�t&}+�QP�������  �jj+�PQ�������  3�3�9M�~w�U���X������<������u.�r�4��2������t��r�������t��r�������t���2�4��r�������t��r�������t���X����A��;M�|��M3�Wj�D�  ���_  ���BH�u��HxWh'  V�у��E�;���  ��l��������;�t,}+�QP��������
  �jj+�PQ�������`  ��l�����8���;�t&}+�QP��$����  �jj+�PQ��$�����  3�3�9uȉ}���  ���$    ����ٕx�����p���ٕt���Qٕp���W�U��U�ٕ|����U��U��U��U��U��]��BD�Uċ@<R�Ћ�X����v�����<���   ��������U���U��Q�U��Q�������U��T�U��D�M��H�P�������F�@����|�����U��Q�U��Q�������N�I����p����:��t����z��x����z��(����4���(����V�T���(����}�����(������   �������U���U��T�U��T��|���ȋ������T�U��D�M��H�P�������F�@����p������t����Q��x����Q��(����4���(����V�T���(�������X���4�G;}ȉ}��M����MȋU��uQ�M�R�U�������PQRV���;���������Cj j����  ��t	�����K�������E�"��������\������   �M苐�   G��\�����;������3��M��@ 9�����t9{~�UVR���������H�Al��D���R�E�!�ЍM�Q�E���? �U�R�}��E���? ���z  j h�t��`����m���3�Vhlt�M��E�3�Y��������   �M��Bx�E�4��P�M�Q������R�a  ��`���QP�������5R�]��H  P�E�6讇 ���H�Al������R�]��Ћ��Q�Jl������P�E�4�ы��B�Pl�M�Q�E�3�ҡ��H�Al��`���R�E�0�Ѓ�,�������E�"�~������Q�Jl��D���P�E�!�эU�R�E���> �u��E�P�E���> ���M�u��E���  �����������E�"�"������Q�Jl��D���P�E�!�эU�R�E��|> �E�P�E�    �E��h> ���E�    ���   ���   �E�P�E��у��E�    �#������B�P`�M�Q�ҡ��H�AdWj��U�h8tR�Ћ��Q�J`�E�P�E�:�ы��B�PdWj��M�h,tQ�҃�(�����   �Bx���E�;��P�M�Q������R�  �M�QP�������<R�]��k  P�E�=�х ���H�Al������R�]��Ћ��Q�Jl������P�E�;�ы��B�Pl�M�Q�E�:���E�0���H�Al�U�R�Ѓ�,�������E�"褰�����Q�Jl��D���P�E�!�эU�R�E���< �E�P�}��E���< ���}싑�   ���   �E�P�E��у��}��������H�A`�����R�Ћ��Q�Jdj j������htP�э����R�E�>� ���H�Al�����R�E��Ѓ�3��� ���Q�)� �����   ���   �M�Q�E��҃��������}��E��X8 �������E� �I8 �������E������78 �   �M�d�    Y_^[��]� �������������̡�V�񋈜   ���   V�҃��    ^���������������V��V�; ���    ^�������������U��Q3�9A~V�u�2@��;A|�^]� ���������������U���VW�}���}
_3�^��]� �F;ǉE����ES�E��]��M���r�������*  )^�F��   �؉E�E���v�]�E�$�O �]�F�M�W FF���P�N�I���  j ��j P�у��E���%  ��~M�N�ۍI�N�S��PQ�~����F�M+Ǎ@�F�E�ҍ@R���FR�P�T����]���!�N�I��Q�N�I�N��PQ�.�����V��V �F�M�@������F�b  ��@���F���O  ���Q�[��QP�R ���2  �VщU�E���v�]�E�$��M �]�F���M��U ��;^�]���   ���H���  �[j ��j R�Ѓ��E��u[_3�^��]� �N;�}M�N�ۍIۍ��FSRP�K����F+Ǎ@�F�Eɍ@�E�Q���VQ�R�!����]�����I��Q�N�I�N��PQ�������V�U �F�M�@������F�^�/�F;�}(�N+Ǎ@��R����E�R�@��P�Q ���]�} tC�N;�} ��+��@��R�I�N��j R�J ���V�[��P���j P�tJ ���} tO�N��;�}!�F�I����+х�t�P�P�����u�V�����~�˅�t�P�P�����u��؋E�[�F_�   ^��]� ��������U��QVW�}����  �N;��M��  �> ��  �E��;�u���$	  _�   ^��]� S�;�|���E+��E���r������A�_  ^�F�N;��E�M�
  �E���]�E�u�]��E��$�^J �]��E��M�S )F�V�M+ȉN���H���  �Rj ��j R�Ѓ��E���H  ��~O���Q�N�I�N��PQ�����F�M+�+Ǎ@�F���R�@���N�R���R躛�����)�N+ˍI��Q�N�I���VP�[��P菛����V�FS �F�M��)^�@[���F_��   ^��]� ��~�F���QP�[��P�O ���F�)^�@[���F_�   ^��]� +�N���M�E�v�]�E�$�DJ �]�F���M�3R ;F�E��   ���Q���  �@j ��j P�у��E��u[_3�^��]� �N�Q�;�}O���Q�N�I�N��PQ萚���F�M+�+Ǎ@�F���R�@���N�R���R�a������ +ˍI��Q�N�I�N��PQ�?�����V��Q �F�M��)^�@����M[�F_�N�   ^��]� �F�P�;�}(�N+�+Ǎ@��P�;�@��P���P�M ��)^[_�   ^��]� _3�^��]� ��������������U���VW�}���}
_3�^��]� �F;ǉE����ES�E��]��M���r�������
  )^�F��   �؉E�E���v�]�E�$�~H �]�F�M�pP FF���N�Pj ��    ���  j P�ы؃����  ��~E�V�N��    P��PQ�����V�F+���E�R�V����    Q�R躘������F�N��P�F��RP蝘����V�TP �N����]���V�3  ����F���#  ��    R��QP�	  �VщU�E���v�]�E�$�}G �]�F���M�lO ;F�E��   ���Q���  j ��j P�ы؃���u[_3�^��]� �F;�}E�V�N��    P��PQ�ӗ���V�F+���E�R�V����    Q�R諗������N��P�F��RP著����V�HO �N�E����]���V�F�$�F;�}�N+���P���R��Q�K ���} t:�F;�}�N��+���R��j R�7D ���N��    P��j R�D ���E�[�F_�   ^��]� �������U��QVW�}�����  �N;��M���  �> ��  �E��;�u���$  _�   ^��]� S�;�|���E+��E���r������A�9  ^�F�N;��E�M��   �E���]�E�u�]��E��$�^D �]��E��M�M )F�M�V+ȉN���H���  j ��j R�Ѓ��E���"  �V����~>��    Q�NPQ�����V�F�M+�+���RǍ��NR�;��R�ȕ������N+���Q�NP��R謕����V�cM �E�N��)^[���_�V�   ^��]� ��~�F��    QP��R�8I ���F�)^[��_�V�   ^��]� +�N���M�E�v�]�E�$�jD �]�F���M�YL ;F�E��   ���Q���  j ��j P�у��E��u[_3�^��]� �N�Q�;�}D�V��    Q�N��PQ輔���V�F�M+�+���RǍ��NR�;��R蕔�����+���Q�N���FRP�y�����V�0L �E�N��)^����E[�F_�V�   ^��]� �F�H�;�}�N+�+���P�;��P��Q��G ��)^[_�   ^��]� _3�^��]� ����U���V��H�QV�ҋ��Q�M�R0QPV�҃���^]� ��������������U����P�Ej PQ�J �у����@]� �������������VW��3�9>t	V�@K ���>�~�~�~�~_^�������������U��Q�E;�u	�   ]� }+�RP�O���]� jj+�PR�~���]� ����������U��j�hAXd�    P��V�p�3�P�E�d�    �E�    ���H�A`�U�R�Ћ��Q�M�Rp�E�PQ�ҡ��H�A�U�R�E�   �Ћ��Q�MQ�J0P�E�P�ы��B�u�H`V�ы��B�Pp�M�VQ�ҡ��H�Al�U�R�E�   �E� �Ѓ�,�ƋM�d�    Y^��]��������U��V��W�~��}_3�^]� jjjW�n�����t�F�M��_�   ^]� �������Du�J �����U��V���Du�J �Et	V�CN ����^]� ���������U��M�UV�uW��r�;u��������s��tE��9+�u1��v6�B�y+�u ��v%�B�y+�u��v�B�I+���_��^]�_3�^]�����������U��QV��j �M��. �F���s@�F�M��. ^��]�������U��QVW��j �M���- �G��v	���sH�G�w����֍M�#���- _��^��]�����Pu����������U��QW�9��t=j �M��}- �G��v	���sH�GV�w����֍M�#��- ��t
��j����^_��]����U���EV���Put	V��L ����^]� �������������̰�������������̸   �����������U��Q�A$V�0W�}j �M�E�    �7��, �F���s@�F�M��, ��_^��]� �U��V��V�Xu�0 ���Et	V�/L ����^]� �����U��j�hyXd�    PQVW�p�3�P�E�d�    ���E�    �u���E�    衽  ���H@�Q`VW�E�    �E�   �҃��ƋM�d�    Y_^��]� �����������̡��P�Bl��Q��Y��������������U��MV3��r� ��t�����   ���ȋB(�Ѕ�u��^]� ��������������U��j�h�Xd�    P��SVW�p�3�P�E�d�    ���E�    �j� �O ���EP��S P���� �M�Q�������jh�  �M��E����  jh�  �M����  �URh�  �M����  jh�  �M����  ���H@�Adj�U�RV�Ћ]����3�脧 ��t�����   ���ȋB(�Ѕ�u�WV����� �����   �Bj j���ЍM��E� 苼  ���Q�Jl�EP�E������у��M�d�    Y_^[��]� �����������U��j�h�Xd�    P��4SVW�p�3�P�E�d�    ��u���HT�U�A,j R�Ѓ��E��u�M�d�    Y_^[��]� �M�Q���� ���   +��   �]�ƨ   ���g������������E�    ;�r�6I �N��i��   �T9Rh�  �M��2�  �N+N���g�����������;�r��H �N��9�    tIS���S  ��LPh�  �M��*�  �U���R�M��[# �E�Ph�  �M��E��&�  �M��E� �# �M�Q�M�n� �M��E��������  �   �M�d�    Y_^[��]� ������U��j�h6Yd�    P��TSVW�p�3�P�E�d�    ���}���H�A`�U�R�Ћ��Q�Jdj j��E�h�rP�у����   +��   �]�Ǩ   ���g������������E�    ;�r��G ���Q�R ��i��   Gj �M�Q��\P�ҋ���H�Al�ލU��R���E������Ѓ�����  ���QT�u�B,j	V��3Ƀ��E;�u3��M�d�    Y_^[��]� �M�M�h�  �M��E�   �^� j �M�QP���E��̘ �M��E�谄 �E�   �E�    �����   �@�M�Q�U�R�E��Ћ����   �
�E�E�P�E��у��} tW�E�   �E�   h�  �M��E��ґ j �U�RP���E��`� �M��E��$� �����   ��U�R�E��Ѓ��u�M�Q���� S���E�� Q  ��4Ph�  �M��_�  S����P  ���    tIS����P  ��\Ph�  �M��u�  �U���R�M��  �E�Ph�  �M��E��q�  �M��E���  �M�Q���� �M��E��N�  �����   ��M�Q�E������҃��   �M�d�    Y_^[��]� �������U��j�h�Yd�    P��TSVW�p�3�P�E�d�    ���}���H�A`�U�R�Ћ��Q�Jd3�Sj��E�h�rP�у����   +��   �u�Ǩ   ���g����������]�;�r�E ���Q�R ��i��   GS�M�Q��pP�ҋ���H�Al�ލU��R���E������Ѓ�;���  ���QT�u�B,jV�Ѓ��E;�u3��M�d�    Y_^[��]� �]�]�h�  �M��E�   蔏 S�M�QP���E��� �M��E��� �E�   �]�����   �@�M�Q�U�R�E��Ћ����   �
�؍E�P�E��у���tW�E�   �E�   �h�  �M؈]��� j �U�RP���E�蝕 �M؈]��b� �����   ��U�R�E��Ѓ��]�M�Q���J� �uV���E��;N  ���    tIV���*N  ��pPh�  �M��ɾ  �U���R�M��� �E�Ph�  �M��E��ž  �M��E��9 �M�Q���� �M��E�袵  �����   ��M�Q�E������҃��   �M�d�    Y_^[��]� �����������U��j�h�Yd�    P��TSVW�p�3�P�E�d�    ���}���H�A`�U�R�Ћ��Q�Jdj j��E�h�rP�у����   +��   �]�Ǩ   ���g������������E�    ;�r�SB ���Q�R ��i��   Gj �M�Q��pP�ҋ���H�Al�ލU��R���E������Ѓ����  ���QT�u�B,jV��3Ƀ��E;�u3��M�d�    Y_^[��]� �M�M�h�  �M��E�   �ތ j �M�QP���E��L� �M��E��0 �E�   �E�    �����   �@�M�Q�U�R�E��Ћ����   �
�E�E�P�E��у��} tW�E�   �E�   h�  �M��E��R� j �U�RP���E���� �M��E��~ �����   ��U�R�E��Ѓ��M�Q�M�� S���K  �@l�5�u�E�   �]�E�]�h  �M��E��܋ j �U�RP���E��j� �M��E��.~ �����   ��U�R�E��Ѓ�S���K  ���    tIS���K  ��pPh�  �M�誻  �M���Q�M��� �U�Rh�  �M��E�	覻  �M��E�� �M�E�P��� �M��E�育  �����   �
�E�P�E������у��   �M�d�    Y_^[��]� �����������U��j�hgZd�    P��TSVW�p�3�P�E�d�    ���}���H�A`�U�R�Ћ��Q�Jdj j��E�h�rP�у����   +��   �u�Ǩ   ���g������������E�    ;�r�3? ���Q�R ��i��   Gj �M�Q��P�ҋ���H�Al�ލU��R���E������Ѓ��   ����  ���QT�u�B,jV��3Ƀ��E;�u3��M�d�    Y_^[��]� �M��M�h�  �M؉]�轉 j �M�QP���E��+� �M؈]��| �E�   �E�    �����   �@�M�Q�U�R�E��Ћ����   �
�E��E�P�]��у��}� tR�E�   �]�h�  �M��E��7� j �U�RP���E��ŏ �M��E��{ �����   ��U�R�]��Ѓ��M�Q�M�t� �E�   �]�h�  �M��E��و j �U�RP���E��g� �M��E��+{ �����   ��U�R�E��Ћu��V���H  ���    tIV���H  ��Ph�  �M�褸  �M��Q�M��� �U�Rh�  �M��E�	蠸  �M��E�� �M�E�P�� �M��]��}�  �����   �
�E�P�E������у��ËM�d�    Y_^[��]� ���������U��j�h�Zd�    P���  �p�3ŉE�SVWP�E�d�    ���V ��ٕH�����T���ٕL�����H���� uPٝP��������Q�����ٕ���R�荅8���ٕ���3�ٝ���P��������X���ٕ ���ٕ���ٕ���ٕ8���ٕ<���ٝ@����~�����Q�J`��4���P�ы��B�PdVj���4���hxvQ�ҍ�4���P�u��c ���Q�Jl��4���P�E������ы��   +��   �����������������\�����
  ��`������   +��   ���������������9�\���r�N; ���   �`����{ �   ��x������   ���B�P`��4���Q�ҡ��H�Idj j���x���R��4���P�у���T�����4���R�E�   �D ��D������H�Al��4���R�E������Ѓ���D��� t��D���Q軧 ���U܋E�RP�� ������h�������	  ���   +��   ���������������9�\���r�S: ���B���   �P`�`��������Q�ҡ��H�Adj j������WR�Ѓ������   �R|�����P���E�   �ҡ��H�Al�����R�E������Ћ��QH�B|j h�  V�Ћ��QHj ��t����B|h�  V�Ѓ��}� ǅp���    ~o3��
��$    �I �U�t��X���+���d����t+���l����t�+׉��l���+��p�P��d����P��p���B�� ��;U܉�p���|���h���3�9}���   ��X���م����م������t���م�����Rم�����م����ҋ��   ��؍����G����؅�����@؍���������H��ٝt���� ؍����؅�����@�������H��ٝl���� ؍����؅�����@�������H��ٝp���مt���ٝH�����H���مl����A�ٝL�����L���مp����A�ٝP�����P����A�;}��>������������؃; ��  �}� ��  ��M�ٕ����Qٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٝ������� ������l������$  �}� ǅp���    �  3���d������d����M�T�t�|���   �<�<���t�����d����L�I�R���4v�4������P����H�@��X�����t�����T������\����H�@��`������d����F��h����N��l������p����J�R��t�������x�����|����   ��P����������HD��p���������R��l���P�A@R�Ћ�p�����d��� @��;E܉�p����������l�����h���j W���4� �����   �Bj j����j h�  ��迓 ����   ���Q�J`�����P�ы��B�Pd3�Wj������hPvQ�҃������   �Bx���E�   ��P�����Q�����R�s���P�E���\ ���H�Al�����R�E��Ћ��Q�Jl�����P�E������у��3�9{��  ���B�P`��$���Q�ҡ��H�AdWj���$���h�rR�Ѓ����   +��   ���g����������ʃ����   �E�   ���g�un+��   ��$���R����������u� 5 ���   ���B����t����H`����l���W�ы��B��t����PpWQ�҃�V��������  +��   ������������  ��$���Q���   +��   ���g�����������u�j4 ���   ���B����t����H`����l���W�ы��B��t����PpWQ�҃�V���������   +��   ���g�����������   �;��?  ǅp����   h)  �̿ ���Q������l������0  �J`��@���P�ы��B�Pdj j���@���hDvQ�ҍ� ���WP�E��%� P��@���Q��0���R�E��������Q�Rp��$���QP�E��ҡ��H�Al��0���R�E��Ћ��Q�Jl�� ���P�E��ы��B�Pl��@���Q�E��ҡ����   �R|��<��$���P���ҋ�覻 3�9u܉�t���~�E�9<�u��t���V�� F;u�|拍h���3��� ��t�����   ���ȋB(�Ѕ�u狍h���V��l���V�R� �����   �Bj j���Ѝ�$���Q���   +��   ���g�����������;�r�C2 ���Q���   �p������ĉ�t�����t���P�B`�Ћ���t����Q�JpPV�ы�h�����R����������   +��   ��p����   ���g����������G�;��������h���3����Q�Jl��$���P�E������у���T���jWWV�7 �����   �PWj���҉������������������������� ���ǅ����   ��������T���������Qh�   �E�	   �������������Y ���E���������������   �U��X����\�  ���   +��   ��\�����`���x��������������F�\���;��>����   �M�d�    Y_^[�M�3��� ��]ËJl��$���P�E������у�3�����  3����������������U��j�h [d�    P��SVW�p�3�P�E�d�    �񋎸   +��   ���g����������3���-  �]����   +��   ���g�����������;�r��/ ���   E��N P��8 ����uihG  �B� ��������   ���   +��   ���g�����������;�r�/ �����   ���   E��R|P���ҋN j j W�S5 WS������WS��������~ W��Su�b��������WS���r���jj���� �����   �Bj j���Ћ��   +��   �E�   ���g����������C�;�������   �M�d�    Y_^[��]Ë��B�P`�M�Q�ҡ��H�Adj j��U�h�vR�ЍM�Q�E�    �U ���B�Pl�M�Q�E������҃�3��M�d�    Y_^[��]����������������U��j�hr[d�    PQSV�p�3�P�E�d�    ��u����   P�E�   �. ���   P�w. �����   �y  ���   3�;�t	P�. �����   P���   ���   ���   ��- ���N\�E�� �N@�E�� �N$�]�� ���H�Ql��V�E������҃��M�d�    Y^[��]�����U��j�h�[d�    P��SVW�p�3�P�E�d�    ��u���Q�FP�B`�Ѓ��N$�E�    �o �N@�E��c �N\�E��W ���   ���E��F�  ���   ���E��5�  3��Fx�F|���   ǆ�   �����G�E��E�9Gv��, ��M��O�M�;Ov�, �M��U�R�U�RQP�E�P����a  �{9{v�, ��M��K�M�;Kv�o, �M�U��WRQP�E�P���o  �ƋM�d�    Y_^[��]��������������U��j�h:\d�    P��\  �p�3ŉE�SVWP�E�d�    �u�ٿ   W��0����\�  j@WV��8����E�    �f�  ��u+��0����H��8�����0������y( u��j P�u  ������ ��  ���Q�J`������P�ы��B�Pdj j�������h�wQ�ҡ��H�A`������R�E��Ћ��Q�Jdj j�������huP�ы��B�P`������Q�E��ҡ��H�Adj j�������VR�Ѝ�����Q������R������P�]�������H������QP�� ���R�E��e���P�E���Q ���H�Al�� ���R�E��Ћ��]��Q�Jl�����P�ы��B�Pl������Q�E��ҡ��H�Al������R�E��Ћ��Q�Jl������P�E� �у�$�������E������܀  ������Rǅ����Xu� ��3��F  ���H�A`������R�Ћ��Q�Jdj j�������h�wP�э�����R�E��Q ���H�Al������R�E� �Ћ�0����A��8��������c  j
��0����(v  ��Rjc������P��0������  j������QhDs�>5 ����uG{|���   +��   ���   ���������������;�r�,) ���   ����+΍D�h��  j������Ph�w��4 ����uJ��   ���   +��   ���   ���������������;�r��( ���   ����+֍D�l�_  j������Qh�s�y4 �����  ��   ���   jx������@j R�������: ��l���   ������󥋍�������   Q���  ���   +��   ���   ���������������;�r�( ���   ����+�3��|�d���   +��   ���   ���������������;�r��' ���   ����+Ή|�h���   +��   ���   ���������������;�r�' ���   ����+Ή|�l�   �4j������Ph�w�L3 ����u���   {xQ���   �1  ��d8��0����B��8����������8����hk  ��u+��0����H��8�����0������y( u��j P�ip  �s|3ɋƺ   �������Q�# �����t�V���|�H�Q�����Q��Q�y��3����   �؉��   3ɋƺ   �������Q�`# ����t!�V���|��H�Q�����Q��Q�y����3����   ���   +��   ��������������3���C  3����   +��   ���������������;�r�& ���   ǋ@d3�@�    �������Q�" ���   +��   ���������������������;�r��% ���   �������Tp���   +��   ���������������;�r�% ���   ǋ@d3�@�   �������Q�2" ���   +��   ���������������������;�r�8% ���   �������T9t���   +��   ��������������F�x;�������������E������{  ������Qǅ����Xu�v	 ���   �M�d�    Y_^[�M�3��� ��]� ��������U��j�h�]d�    P��l  �p�3ŉE�SVWP�E�d�    ��j�������ӄ  �������^\P���E�    �  ���Q�JP������jP�E��ы����B��H  j Gj W�ы��JjWP�������������ATR�Ћ�������$j@jQ�������o}  ��u+�������J���������������y( u��j P� m  ������ ��  ���H�A`��p���R�Ћ��Q�Jdj j���p���h�wP�ы��B�P`��`���Q�E��ҡ��H�Adj j���`���huR�Ѓ�(��(���Q���E����  P��`���R�� ���P�E�������p���QP������R�]�����P�E���I ���H�Al�����R�]��Ћ��Q�Jl�� ���P�E��ы��B�Pl��(���Q�E��ҡ��H�Al��`���R�E��Ћ��Q�Jl��p���P�E��ы��B�Pl������Q�E� �҃�4�� ����E�������x  �� ���Pǅ ���Xu�� ��3��b  ���Q�J`��`���P�ы��B�Pdj j���`���h�xQ�ҡ��H�A`��p���R�E��Ћ��Q�Jdj j���p���huP�у�(�����R���E��u�  P��p���P�� ���Q�E�	�-�����`���RP��(���P�E�
����P�E��{H ���Q�Jl��(���P�E�
�ы��B�Pl�� ���Q�E�	�ҡ��H�Al�����R�E����E����Q�Jl��p���P�ы��B�Pl��`���Q�E��ҋ������@��������0�������  �l����������	�I ������j
�������Lm  ��Qh�   ������R��������  j������Pht�_, �����  ��   �Ô   ��G��������������+  �O���   Q���x  ������R������h�xP�e- ���Q�J`��p���P�ы��B�@dj j�������Q��p���R�Ѓ� �K+K���g������������E�;�r�� �C��������JP�Ap��p���R�Ћ��Q�Jl��p���P�E��ыK+K���g�����������;�r�v �K������Ǆ
�       ��  j������Ph�x�$+ ����������u^�����Qh�xR�_, ���   +��   ���g�����������;�r�  ݅������   ٝ����م�����\�q  jRh�x�* ����ud�����P������h�xQ��+ ���   +��   ���g�����������;�r� ݅������   ٝ����م�����\��  j������Rh�x�.* ����u)W���   ��(  ��P������h�xP�`+ ���  j������Qh�x��) ������   ��X���R��H���P��P���Q������hxxR�+ ݅P�����ٝ�������   W���l(  م�����XW݅H�����ٝ�����O(  م����W�X ��݅X���ٝ�����2(  م�����X$�  j������Phtx�B) ������   ��X���Q��H���R��P���P������hdxQ�k* ݅P�����ٝ�������   W����'  م�����X(W݅H�����ٝ�����'  م����W�X,��݅X���ٝ�����'  م�����X0�d  j������Rh`x�( ������   ��X���P��H���Q��P���R������hPxP��) ݅P�����ٝ�������   W���'  م�����X4W݅H�����ٝ������&  م����W�X8��݅X���ٝ������&  م�����X<�  j������QhLx��' ������   ��X���R��H���P��P���Q������h<xR�) ݅P�����ٝ�������   W���q&  م�����X@W݅H�����ٝ�����T&  م����W�XD��݅X���ٝ�����7&  م�����XH�  j������Ph4x�G' ����uZ������Q������h(xR�( ��j ������P�������J��������Q���   W���E���%  �ȃ�L�\���������vj������Ph x��& ������   ������Q������hxR�
( ��j ������P�������(J��������Q���   W���E��O%  �ȃ�\�\�����������B�PlQ�E��҃�W���!%  ǀ�      �������@������������������^  ��u+�������I���������������y( u��j P�c  j��D����yz  ��4����^@R���E����  ���H�AP��4���jR�E��Ћ��Q����H  j Gj W�Ћ��Q�JTjWP��������4���P�ы�������$j@jR��L����s  ��u+��D����H��L�����D������y( u��j P��b  ������ ���Q�J`��`���P��  �ы��B�Pdj j���`���h�wQ�ҡ��H�A`��p���R�E��Ћ��Q�Jdj j���p���huP�у�(�����R���E���  P��p���P�� ���Q�E��W�����`���RP��(����P�]��>���P�E��? ���Q�Jl��(���P�]��ы��B�Pl�� ���Q�E��ҡ��H�Al�����R�E��Ћ��Q��p����E�P�Jl�ы��B�Pl��`���Q�E��ҡ��H�Al��4���R�E��Ѓ�4�������E��n  �������XuQ�������� ���B�Pl������Q�E� �҃��� ����E������Zn  �� ���P�� ����@� ��3���  �ы��B�Pdj j���`���h�xQ�ҡ��H�A`��p���R�E��Ћ��Q�Jdj j���p���huP�у�(�����R���E����  P��p���P�� ���Q�E�������`���RP��(����P�]�����P�E���= ���Q�Jl��(���P�]��ы��B�Pl�� ���Q�E��ҡ��H�Al�����R�E��Ћ��Q��p����E�P�Jl�ы��B�Pl��`���Q�E��ҋ�D����@3���0��L�����������  j
��D�����b  ��Qh�   ������R��D����rx  ���   +��   ���g����������3����   ���������Q�J`��p���P�ы��B�@dj j�������Q��p���R�Ѓ����   +��   ���g������������E�;�r� ���J���   �����j ��p���RP�A �Ћ��Q�Jl���ߍ�p����PG�E��у���u4���   +��   �������   ���g����������C�;������������������j������Qhx��  �����*  ���   +��   ���g�����������;�r�� ���   i��   �TlR������h�wP��! ��D����I��j
��D����$a  ��Rh�   ������P��D����v  ���Q�J`��`���P�ы��B�@dj j�������Q��`���R�Ѓ����   +��   ���g������������E�9�����r� ���   ���H�Ap�|p��`���WR�Ћ��Q�Jl��`���P�E��ы�������   j	������Rh�w� ������   ��D����Hj
��D����)`  ��Qh�   ������R��D����u  ���H�A`��8���R�Ћ��Q�Rdj j�������P��8���Q�҃����   +��   ���g������������E�;�r� ���   ��iɔ   ���   ���Q�JpP��8���P�ы��B�Pl��8���Q�E��҃���D����@��L����b���3���L���9�����t ���fH  ��u3�������Q�� ����t3���T�����\�����X�����d�����h�����`�����l�����p�������t�����x���ƅ���� ƅ���� ��|�����������X�����h�����x�����T�����d�����t���������������������;�u)��D����H��L�����D�����9y(u��WP�,[  ������V�Q ������Y  ���Q�J`������P�ы��B�PdWj�������h�wQ�ҡ��H�A`������R�E��Ћ��Q�JdWj�������huP�ы��B�P`��8���Q�E��ҡ��H�AdWj���8���VR�Ѝ�8���Q������R������P�E� ������H������QP�������!R�]��r���P�E�"��7 ���H�Al������R�]��Ћ��E� �Q�Jl������P�ы��B�Pl��8���Q�E��ҡ��H�Al������R�E��Ћ��Q�Jl������P�E��у�$���B�Pl��4���Q�E��҃��������E���f  �������XuP�������� ���Q�Jl������P�E� �у��� ����E������f  �� ���R�� ����q� ���   �M�d�    Y_^[�M�3���� ��]������V����������1����   ^�����������U��j�h4^d�    P��$SVW�p�3�P�E�d�    3��u�M�u��e  �E�]jV�M�Q�ˉu��E�   �E���)  �������   �U�U��    ��+�PV�M�Q���L  �MP�E�   �_{  �}��E� r�U�R� ��j�wV�EP���)  �����u�PV�M�Q���4L  �uP���E�   �{  �}�r�U�R�� ���ƋM�d�    Y_^[��]� �E�M�d�    Y_^[��]� ���U��j�hm_d�    P��  �p�3ŉE�SVWP�E�d�    �]����������������@����fd  3��������u��Vd  j�������E��en  j@jS�������E��qg  ��u)�������H��������������9q(u��VP�$W  9�������  ���Q�J`��d���P�ы��B�PdVj���d���h�wQ�ҡ��H�A`��T���R�E��Ћ��Q�JdVj���T���huP�ы��B�P`������Q�E��ҡ��H�AdVj�������SR�Ѝ�����Q��T���R��(���P�E�蒽����H��d���QP��D����R�]��v���P�E���3 ���H�Al��D���R�]��Ћ��E��Q�Jl��(���P�ы��B�Pl������Q�E��ҡ��H�Al��T���R�E��Ћ��Q�Jl��d���P�E��у�$�������E���b  ������Rǅ����Xu��� ���������Lh  �������Ah  3��  ���H�A`��d���R�Ћ��Q�JdVj���d���h(yP�ы��B�P`��T���Q�E��ҡ��H�AdVj���T���hyR�Ћ��Q�J`������P�E�	�ы��B�PdVj�������SQ�ҍ�����P��T���Q��(���R�E�
�������H��d���QP��D����R�]��ػ��P�E��>2 ���H�Al��D���R�]��Ћ��E�
�Q�Jl��(���P�ы��B�Pl������Q�E�	�ҡ��H�Al��T���R�E��Ћ��Q�Jl��d���P�E��ы��B�P`��l������Q�������������ҡ��H�A`������R�E��������Ћ��Q�JdVS������hyP�э�����R�E��&2 ���H�Al��������@R�E��Ћ������A������������	  3ۉ������������j
�������V  ��Rh�   ������P�������'l  j������Qh�s� ������   ������R������h yP�� ��@�����Q��t������  ��t����w\R���E��g�  ��t����E��h�  ����  ������P��t�����  ��t���Q���E���  ��t����E��.�  ��  j������Rh�s�� ������  ���H�A`������R�Ѓ��������������E���;�v�� ��������������������;�v�� ������SVWQ��\���R�������g  �   3�������������������ƅx��� �P�@��u�+�P������P��t����9  jj��t���Q��l����E��i  �   9�����r��x���R�^ ��������P�� �ĉ8�p�x������������ƅx��� �������@ �� ��l����̉�����R�E���r  ������P�E���u  ������������+θ�$I����������ʃ�H��w� ������9^4r�v ��� ���B�P`��D���Q�ҡ��H�AdWj���D���VR�Ћ��Q�Rp������P��D���Q�E��ҡ��H�Al��D���R�E��Ћ��������   +��   �ƨ   ���g������������ �tw3ۍ�$    �N+N���g�����������;�r�� ���Q�F�R j �������QP�҃����   �N+N���g����������GÔ   ;�r��N+N���g������������   �|
�̉�������  W���^  �N+N���g���ыN+N������x����g�����������;�r� ��i��   ~�Q�Jp������WP�ыN+N���g�����������L��������������E��\'  ������Rǅ����Xu�N� ���H�Al������R�E��Ѓ��*  �������j������Qh�s�L ����u9������@P���   �������������  P������h�xR�n ����  j������PhDs�� ������   ��0���Q��|���R������P������h�xQ�" ݅����������ٝ�������   م��������   ݅|�����ٝ������م�����\����   ݅0���ٝ����م�����������\��/  j������Ph�w�K ������   ��8���Q�� ���R������h�xP�{ ��l���Q��8���R�� ���P������h�xQ�U ݅ ������   ٝ����م������$����   ���ܥ8���ٝ����م�����\����   ݅l���ٝ����م�����������\��f  j������Rh�w� �����H  ���������t������P���   ��  �Ht���������������c  ������P��P����@  jj��P���Q��l����E��d  ��P����-  ������R�� �ĉ0�@   �p�������@ �� ��l����̉�����P�E��n  ������Q�E���p  ��H��������b  ��������������+˸�$I�����������   �;��L  �����������   ��������$    ������j/V�������\  P��x���R�������P�������E��mh  ��x����E��n^  j �������!  �xr�@���P�z �X����������ǐ   P���s  �Hp�������\�j��������  �Hj h�rQj ���U  ��tJj�������  �xr�@���P� ��������R�ύX��  �������@p���Ή\���������������������+˸�$I����������F�;������+���$I�������������   j �������  �xr�@���P�r ���������������������ǐ   Q�ύX����\  �Pph�rj�������\2��  P�,  ����t<j�������  �xr�@���P� �X���������P���  �Hp�\1�������������E��"  ������Rǅ����Xu�� ��������������3��������@�������7���������9�����t ����5  ��u3�������Q�u ����t3���������������������������������������������������������������ƅ���� ƅ���� ������������������������������������������������������������������;�u)�������H��������������9q(u��VP�H  ���Q�Jl��l���P�E��у��������E���U  ������Rǅ����Xu�� ��������;�t*������Q������������RQP�G  ������R��  ��������P���������������������  ��������;�t*������Q������������RQP�F  ������R��  ��������P��������������������  ���   �M�d�    Y_^[�M�3��i� ��]� �������U��j�h�`d�    P��<  �p�3ŉE�SVWP�E�d�    �}�E��j j	�ωF ��r  j j�ω��r  j j�ωF��r  j j
�ωF�s  �F���Q�J`������P�у�������Rj������P���E�    �*u  ���R�NQP�Bp�E��Ћ��Q�Jl������P�E� �ы��B�Pl������Q�E������ҡ��H�A`������R�Ѓ�������Qj������R���E�   �t  �E�P��������  �������^$P���E���  �������E����  ���Q�Jl������P�E��ы��B�Pl������Q�E������҃�hDr���������  ������P���E�   �H�  �������E������f�  ���Q�J`������P�у�������Rj������P���E�   ��s  P�������E����  �������~@Q���E���  �������E����  ���B�Pl������Q�E��ҡ��H�E������Al������R�Ѓ�h,y�������%�  ������Q���E�	   �p�  ����������}���  j��������[  ������R���E�
   �=�  ���Q�RTj h�   ������QP�E��ҡ��H�Al������R�E�
�Ѓ�j@j������Q�������T  ��u+�������J���������������y( u��j P�\D  ����� ���H�A`�V  ������R�Ћ��Q�Jdj W������h�wP�ы��B�P`������Q�E��ҡ��H�Adj W������huR�Ѓ�(������Q���E��4�  P������R������P�E�����������QP��d����R�]��Ӫ��P�E��9! ���H�Al��d���R�]��Ћ��Q�Jl������P�E��ы��B�Pl������Q�E��ҡ��H�E��Al������R�Ћ��Q�Jl������P�E�
�у�0������}��NP  �����Rǅ���Xu�0� ��3��  ������R�Ћ��Q�Jdj W������h(yP�ы��B�P`������Q�E��ҡ��H�Adj W������hyR�Ѓ�(��d���Q���E����  P������R������P�E�薩��������QP�������R�]��}���P�E��� ���H�Al������R�]��Ћ��Q�Jl������P�E��ы��B�Pl��d���Q�E��ҡ��H�E��Al������R�Ћ��Q�Jl������P�E�
�ы������J��0j
��������D  ��Ph�   ������Q�������tZ  �������Y<  ��u+�������J���������������y( u��j P�ZA  ������P� ��;��`  ���Q�J`������P�ы��B�Pdj W������h�wQ�ҡ��H�A`��t���R�E��Ћ��Q�Jdj W��t���huP�ы��B�P`������Q�E��ҡ��H�Idj W������R������P�э�����R��t���P��T���Q�E�跧����H������RP��D����P�]�蛧��P�E�� ���Q�Jl��D���P�]����E����B�Pl��T���Q�ҡ��H�Al������R�E��Ћ��Q�Jl��t���P�E��ы��B�Pl������Q�E�
�҃�$� ������P���0���������Q��������~ t/���   +��   ���g�����������t���������������V���� j h  �e ��������}��L  �����Qǅ���Xu�� ���   �M�d�    Y_^[�M�3���� ��]� ��������Q�Xu�L� Y��̋A��P�D
�`u��U��V��N+N��������������W�}�;�r�k� �V����+�_��^]� �U��V��N+N���g����������W�}�;�r�+� ��i��   F_^]� ���U��V��N+N��$I����������W�}�;�r��� �V��    +�_��^]� ���������������U��V��赧���Et	V���  ����^]� ���������������U��j�had�    PQV�p�3�P�E�d�    ��u���H�Q`V�����V$�FL�V P�V�E�    �V0�V,�V(�V<�V8�V4�VH�VD�^@���Q�B`�Ћ��Q�F\P�B`�E��Ћ��Q�FpP�B`�E��Ћ��Q�J`���   P�E��у��ƋM�d�    Y^��]�U��j�had�    PQV�p�3�P�E�d�    ��u���H�Al���   R�E�   �Ћ��Q�Jl�FpP�E��ы��B�Pl�N\Q�E��ҡ��H�Al�VLR�E� �Ћ��Q�BlV�E������Ѓ��M�d�    Y^��]���U��A�U��Q �E��U+ЋA0�]� ��������������̋A �8 t�I0��3�����������������U��A�U��Q$�E��U+ЋA4�]� ���������������V���F@t�F�Q��  ���V�    �F �     �N0�    �V�    �F$�     �N4�    �f@��F<    ^�������U��Q�A8V�0W�}j �M�E�    �7�� �F���s@�F�M�� ��_^��]� ̍Q�Q �Q�Q$�A�A�Q(�Q0�A�A�Q,�Q4�     �A$�     �Q4�    �A�     �Q �    �A0�     ���������U��j�hiad�    PQSVW�p�3�P�E�d�    ��u���H�Q`V�ҡ��H�}�QpVW���G�^�^L�GS�^�G�F�O�N�W �V �G$�F$�O(�N(�W,�V,�G0�F0�O4�N4�W8�V8�G<�F<�O@�N@�WD�VD�GH�FH���Q�B`�E�    �Ћ��Q�Jp�GLSP�ы��B�H`�^\S�E��ы��B�Pp�O\SQ���Gl�^l���H�Q`�^p�E�S�ҡ��H�Ap�WpSR�Ћ��Q�B`���   S�E��Ћ��Q�Jp���   SP�ы��   ��<���   �ƋM�d�    Y_^[��]� �����U��VW�����u�� ���t��3ҋE����+��G����;Bw��t�	�3�;As��� w��_^]� ���������U��VW�����u�� ���t��3ҋE�4�    +��G���;Bw��t�	�3�;As�k� w��_^]� ���������U��M����w3ɋ���+����R�~�  ����]Ã��3����xsڍEP�M��E    ��� h���M�Q�E�Du�
� ���U��M����w3�iɔ   Q�%�  ����]Ã��3���=�   sߍEP�M��E    �i� h���M�Q�E�Du�� ��������U��M����w3ɍ�    +���R��  ����]Ã��3����sڍEP�M��E    �� h���M�Q�E�Du�J� ���U��EVP���0� �Du��^]� ����U���VW�}��H�QpVW���G�^�G�^�G�F�O�N�W �V �G$�F$�O(�N(�W,�V,�G0�F0�O4�N4�W8�V8�G<�F<�O@�N@�WD�VD�GH�FH���Q�Rp�FLP�OLQ�ҡ��H�Ip�V\R�G\P���Gl�^l���B�@p�NpQ�WpR�Ћ��Q�Rp���   P���   Q�ҋ��   ��(���   _��^]� ���U��S�]V�u;�t#W�}V��������Ɣ   �ǔ   ;�u��_^[]ËE^[]��������U��S�]V�u;�t#W�}��   ��   V������;�u��_^[]ËE^[]��������U��E��V��M�Q�F�pu�Z� ��V�H�N�P�V�@�F����^��]� ���������������U���E��QP�
� ��]� ��������U��S�]V�u;�tW�y�WP��� �F��;�u�_��^[]� U���E��QP�� ��]� ��������U��S�]V�u;�tW�y�WP��� �F��;�u�_��^[]� U��E]� ������U��E�UV�1W��+�W�}WP�FR��_^]� �������������U��S�]VW�}��+�9us�]� �E�MVSPQ�d� ����_^[]� �����������U��E]� ������U��E�UV�1W��+�W�}W�}WP�F(R��_^]� ���������U��S�]VW�}��+�9us��� �E�MVSPQ��� ����_^[]� �����������U��V��F�pu��~�FP��� �}�NQ���  ���E�Put	V��  ����^]� �������̋��Q�D(��t�H�g� ���������V��W�~8��u��t���(���W�R�  ��_�N^�� ����̃��� ���������̃���������������U��U��@R�Uj�R��]� �������̋�� �����������3���������������� ������������̋A$�8 t�I4��3�����������������V���P�҃��u�^ËF0��F ��Q��^����������U��E�X{�3ɉH�H�H]� ���U��E�X{�3ɉH�H�H]�  ���U��A � ��t<�Q;v5�U���t:P�t�A@u"�A0� �A ����t�A ����]� 3�]� ���]� ̋Q V�2��u���^�SW�y0����;�s�_[^��A@u/�A$� ��t&;�w9q<v9A<s�A<��A<+�I ��_[^�_[���^����������������U��SV�q$�W��t9A<s�A<�]����   �A �����   �E��u�A�y<+8�u��'��u��u�A�u��+8����t�5X{��u����   �A� �y<+�;���   +Q0�)�Q ����   �Q$�����   �Q4�ЋA R��AR�R������p��te���t_�E�=X{��u�A�Y<+�u����u�A�u��+��	����u�u��|�A� �Y<+�;�+Q4�)�I$�
����5X{�E_3ɉ0^�H�H�H[]� ��U��E�UVW�y$�4���t9A<s�A<�X{;���   S�]$��tR�Q ���tI��|w�A� �y<+�;�d+Q0�)�Q ��tX�Q$���tO�Q4�ЋA R��AR�R�����4��t-�?��t'��|#�A� �Q<+�;��Q4+��)�I$��X{��[�E3�_�0�H�H�H^]�  ��������������U��V�q���Q�F�D�`uP� Xu�� ���Et	V��  ����^]� ����U��V��W�~8��u��t���Ř��W���  ���N�� �Et	V���  ��_��^]� �������������U��V��W��u������~8��u��t���j���W��  ���N�W� �Et	V�}�  ��_��^]� ��U��Q�U�E�M���u	;A��   SVW�y;�st+�;�wn�   +���yr
���M�	����M��E�WQS�� ������t5�U�ERPV�ϖ������t,�M�+ލ|�WR�^S�Q� ������u�_^���[��]� �E��x�Mr�	_��^+�[��]� �U��SV�uW��9ws�+� �G+Ƌu;�s���]��;�r�Ãr�����MP�EP�W�4�������u;�s
_^���[]� 3�;���_^[]� �U��M����w3�Q�K�  ����]� ���3����s�EP�M��E    �� h���M�Q�E�Du��� ��������������V�����t(��u�� ��xr�H��H�@�9Fr�� �F^����������U��E��u&�yr�I�E�U�]� �E�U���]� �yr�I����UP�EP�Q��� ��]� ���������U��j�h�ad�    P��SVW�p�3�P�E�d�    �ى]�K��u�� j�E�    ��  ������t.��� �� � j �M����8� �G���s@�G�M��L� �3��ˉs8�����ËM�d�    Y_^[��]�U��S�]V�uW���    ��t)��t%�V�F��r����;�w��r� �N�;�v�1� �7�_��_^[]� ������������U��E�M�UV�uPQRV�� ����^]����������������U��E�M�U ��E��   ]� ����U��E�M��   ]� ������������U��E+E�M;�s��]� ����������U��S�]V�u��+θ����������������+ȋE�ȉM��;�t#+�W��I �<���x�   �;�u�E_^[]�^��[]����������������U��S�]V�u��+˸����������������+���ɋыM��+�;�t+�W�M��M��x�<�   ���;�u�_^[]����������������U����US�]V�uW�}2��E��M��E��E�PQRWVS����+��g�����������iɔ   ����_^+�[��]��������U��U�ES�];�tVW��t�   �����x��x;�u�_^[]����������������V��F � ��t=�N0�	��~�F0��F � �V �� ^Å�t�N0�9 ~����F ��Q���	��P���҃��u�^ËF �8 t�N0�9 ~��^Ë�P��^������U��QV3�9uW���u�~nS�]��������~6�M;ȋ�}��G ��UVQRS�`� �G0)0u�)u�G ރ�0�u����P���҃��tF�C�M�u��} �[_��^��]� _��^��]� ������U��QV3�9uW���u�~mS�]���3�����~3�M;ȋ�}��VSP�G$�Q��� �G4)0u�)u�G$ރ�0�u����P�B���Ѓ��tFC�M�u��} �[_��^��]� _��^��]� �������U��j�h�ad�    PQVW�p�3�P�E�d�    �M��A��P�D
��v�q����E�    ��u�����~8��u��t�������W�)�  ���N��� �F��H�D1�`u�M�d�    Y_^��]����������������U���V���F@Wt �~$���t�N<;�s�F4� +��N4��E���u
_3�^��]� �V$�:S��t$�N4����;�s�	�v$�[�Q�_�^��]� �F@u=��u3���F4�N�+ߋ���� s�    ���v������+�;�s��u��u[_���^��]� �P�ND�E���������F��M���vSQ�M�QW������M�����u"�V�~<�:�F$�8�V4�E���F@u7�GPW�V�F$��+�V<� �V��+�+��V$ǉ��+�U��F4��F@t�V�:�F �     �V0�:��F$��F BR�+��RW���?����M��F@t	Q�p�  ���F4�N@��v$��A��E[_�^��]� �����������̋P�8�  Y�������U��S�]V��W9^s�� �F�}+�;�s����v^�N��r�V��V�U��r�V��V+�P�E��P+�Q�R��� �F+ǃ��~�Fr�N_� ��^[]� �N� _��^[]� ��U��} VW�}��t'�~r!�FS���vWSjP�c� ��S�m�  ��[�~�F   �D> _^]� ����U��E�MPQ�� 3҃������]�V��~L t#��Pj��҃��t�FLP��� ����}���^�3�^�U��A � S�]��t,�Q9s%���t�@�;�u�A0� �I �	��@���#�[]� �AL��t$���t�y< u��PQ�j� �����t��[]� ���[]� �V��F ���t�Ћ�V0��;�s�^Ë�PW���ҋ����u_�^Ë�PW���ҋ�_^������������U��V��NLW��tl�U�}��u	��u�G�3�WPRQ�.� ����uG�~L���FH�FA�������t�G�F�F�G�~ �~$�F0�F4�~L���FD_�F<    ��^]� _3�^]� ��������������U��ES�]V���F<    �F@����   ��<tzWS�ND�@������ESPSW�_� ���F@��F<u�N�9�V �:�N0��N@��u7��u�ǋV�:�N$���+ЋF4Ӊ�N �9 u�V�:�F �     �N0�9�N@_^[]� ����������U��V�1W�y��u��� 3��Miɔ   �;xw��t�����3�;xs�� �E�x_�0^]� �����U��j�h�ad�    P��SVW�p�3�P�E�d�    �e����}�E�������v���"�_������������;�s�����+�;�w�4�NQ���E�    ������E�&�E�M�E�@�e�P�E�������E��Ë}�u�]��v �r�G��GSP�E�VRP��� ���r�OQ���  ���M�G�  ��w�_��r��� �M�d�    Y_^[��]� �u�~r�VR��  ��j �F   �F    j �F �^� �������U����US�]V�uW�}2��E��M��E��E�PQRWVS�����+��g�����������i��   ���_^[��]������������U��E�U;�tS�]VW����x�   ���;�u�_^[]�������U��V�uW�};�tS�]S�������Ɣ   ;�u�[_^]�������U��U��v#�ES�]VW��t�   ����J��x��w�_^[]��U��j�h!bd�    P��SVW�p�3�P�E�d�    �e��u�}3ۉu�]���$    ;}tU�u�u��E�;�tW���e����Ɣ   �]��u�ǔ   �ыu�};�t��$    ���	����Ɣ   ;�u�3�SS��� �ƋM�d�    Y_^[��]���V�qP���5���V�Xu�1� ��^�����V��~r�FP��  ��3��F   �F�F^�����������U��VW�y��wP�������V�Xu�ڹ ���Et	W�S�  ����_^]� ��������U��yr�AV�uQP��������^]� V�u�AQP���p�����^]� ���������U��j�hHbd�    PQV�p�3�P�E�d�    ��u������E3ɉM���u�u�   �u���t���t���E�x�Pr�@���QRP��������ƋM�d�    Y^��]� ����U��U��V�p�d$ �@��u��M+�P�ARPj ���������^]���������������U��Q�M�U�E� �E�P�EQ�MR�UPQR���������]�����U��Q�M�U�E� �E�P�EQ�MR�UPQR��������]�����U��j�h�bd�    P��SVW�p�3�P�E�d�    �e��u�}3ۉu�]���$    ;�vL�u�u��E�;�t�EP������O�Ɣ   �]��u�ԋu�};�t���c����Ɣ   ;�u�3�SS�'� �M�d�    Y_^[��]���������������U��V����v�~$r�FP��  ��3��F$   �F �ΈF�(� �Et	V���  ����^]� �����̃y$r�AÍA���U��j�h�bd�    PQSV�p�3�P�E�d�    ��u�3�S�� �   �F�^�]��^�F8�^4�^$�FT�^P�^@�Fp�^l�^\�EPV�E���� ���ƋM�d�    Y^[��]� ������������U��j�h$cd�    PQSVW�p�3�P�E�d�    ��u�V�E�   �9� ���~pr�F\P���  ��3ۿ   �~p�^l�^\�~Tr�F@P���  ���~T�^P�^@�~8r�F$P��  ���~8�^4�^$�~r�FP��  ���~�^�Έ^�E�������� �M�d�    Y_^[��]���V��~r�FP�N�  ��3��F   �F�F^�����������U��S�]V�����+F;�w�o� ����   W�~����v�W� �F;�s9�NQW���<�����vZ�U�FRSP���8����~�~r:�F�8 _��^[]� ��uщ~��r�F_�  ��^[]� �F_�  ��^[]� �F�8 _��^[]� �����U��S�]VW�}��9_s��� ��E+�;�s���M;�uj��W������Sj ������_��^[]� ���v肶 �M�F;�s�FPW���d����M��vj�yr/�I�-��u�~��r�F_�  ��^[]� �F_�  ��^[]� ���~�^r���ËUW�Q�NQP�� ���~�~r��; _��^[]� ����������U��USVW���tF�~�F��r����;�r1��r���ȋ^�;�v��r� �MQ+�RV�������_^[]� �}���v膵 �F;�s�VRW���k�����vY�N�^��r.��,��u�~��r�F_�  ��^[]� �F_�  ��^[]� �ËUWRQP�� ���~�~r��; _��^[]� �����U��Q�UV�uW�}�E� �E�P�ER��QPVW������΃���+΍�_^��]� ����U��V3���j��F�F   P�F�EP�������^]� ��������U��j�hHcd�    P��D�p�3ŉE�SVWP�E�d�    �A � 3҉M�;�t'�A �q0� �6�;�s�A0��A ��Q���K  �AL;��=  9Q<uP�� ������&  ���!  �E�   �U�U�P�U��a� �������  Pj�M��Y����}�E؃��5  ���u̅�t!�ȃ�s�M�;�w�ȃ�s�M؋U��;�v�"� �}�U�E؍Mԃ��t�ȃ�s�M��;�r��� �}�U�E؋ڃ���   ����t�ȃ�s�M�;�w�ȃ�s�M��;�v�� �}�U�E؍Mԃ��t��s�E��;�r�� �}ċO<��R�E�P�E�P�E�P�E�P�E��PV�GDP�҅���   ��~_����   �}���   j�U�R�M��.���������P�E�jP�H� �uӃ��M��������   �M؉M̋�������u��%����E�9E���   �U�E؃���   ����t!�ȃ�s�M�;�w�ȃ�s�M؋]��;�v��� �U�E؍Mԃ��t��s�E؋U��;�r�� �E�+�Pj �M������OLQ�m� ����������M����������M�d�    Y_^[�M�3��y� ��]Íu��b����}�M�Q�M��"������{���+}ȋ����~�UċBL�M��T�NPR��� ������uӍM��w���������U��V�u��W�x�I �@��u�+�PV�p���_^]� ����������U��SVW�}���    ��t�E9Fw;Fv�� �E�]���G9^w;^v�� �]����t;�t�p� �O;�t!�F�E �UR�UR�URQPS��������F��_^[]� ��������U��j�hxcd�    P��,�p�3ŉE�SVWP�E�d�    �y< �M���  �yA ��  ��Pj��҃���m  �   3��E� �M�E؉E��E�   ��s�E��@ �E�    �E؋U����    ����   �؉]̅�t!�ȃ�s�M�;�w�ȃ�s�M؋u��;�v�o� �U�E؍Mԃ��t�ȃ�s�M؋u��;�r�I� �U�E؋}����   ����t$�ȃ�s�M�;�w�ȃ�s�M؋]�ˋ]�;�v�� �U�E؍Mԃ��t��s�E؋U��;�r��� �EЋH<��R�E�P�E��SV��DP�҃� t)��t+���M��7  �>  �]؉]������u��i����E��@A �U�E؃���   ����t!�ȃ�s�M�;�w�ȃ�s�M؋}��;�v�X� �U�E؍Mԃ��t�ȃ�s�M؋}��;�r�2� �U�E؋}�+�tv����   ����t!�ȃ�s�M�;�w�ȃ�s�M؋]��;�v��� �U�E؍Mԃ��t��s�E؋U��;�r��� �EЋHLQWjV�_� ��;�u7�U�E؋MЀyA t4�������Wj�M�����������u������u��h����M������2��
�M��������M�d�    Y_^[�M�3��u� ��]������U��V�uW�};�t����i����Ɣ   ;�u�_^]� ���������U��Q�UV�uW�}�E� �E�P�ER��QPVW�I�����i��   ���_^��]� ����U��Q�U�E� �E�P�ER�U��Q�MPQR�k�������]� ��U��V�u�~r�FP��  ��3��F   �F�F^]� ���U��S�]V�u;�t!W�}j�j V����������;�u��_^[]ËE^[]����������U����p�3ŉE����M;�tT�PS�XV�p�]��YW�x�X�Y�X�Y�X�Y�X�Q�U��q�q�y�Q�P�p�q�Q�P_�p^�Q[�M�3��� ��]� ���U��j�h�cd�    PQV�p�3�P�E�d�    ��u��-� 3��N��vj��A�A   P�E��A�EP�����ƋM�d�    Y^��]� �������U��EVP�������w��^]� ����V����v�~$r�FP�8�  ��3��F$   �F �F��^�Z� ��������������U��j�h�cd�    PQV�p�3�P�E�d�    ��u��]� 3��N�wj��A�A   P�E��A�EP�;����ƋM�d�    Y^��]� �������U��Q�V�u3�j���R�F   �VP�ΉU��V�������^��]� �������������U��j�h�cd�    P��   SVW�p�3�P�E�d�    3ۉ]��}����   9��   j�6�  �����u3��E�;�t2�M�E�P�Y���P��`����E��E�   �"���j P�λ   �����E�   ���t�����`����]�������t�}�r�M�Q��  ���   �M�d�    Y_^[��]�������V���w�~$r�FP�h�  ��3��F$   �F �F��^銿 ��������������U��V���w�~$r�FP�%�  ��3��F$   �F �ΈF�H� �Et	V� �  ����^]� ������U��UV���W�F   �F    �F �x�@��u�+�PR���-���_��^]� �����U��Q�UV�u3��F�F   �E��F�EPRQ��������^��]� �������������V��F��t	P�`�  ���P�F    �F    �F    �@�  ��^������������U��j�h(dd�    P��4�p�3ŉE�SVWP�E�d�    �]�щUЃ��u3��  �B$���t �B4�0�;�s��B$��Q������  �BL����  �z< uP��P�r� �������  ����  �   3��E� �]̉M�E؉E��E�   ��s�E��@ �E�    �E؋U�I ���	  �؉]ȅ�t!�ȃ�s�M�;�w�ȃ�s�M؋u��;�v��� �U�E؍Mԃ��t�ȃ�s�M؋u��;�r��� �U�E؋}����  ����t$�ȃ�s�M�;�w�ȃ�s�M؋]�ˋ]�;�v�� �U�E؍Mԃ��t��s�E؋U��;�r�t� �EЋH<��R�E�P�SV�E�P�E�P�E�P�EЃ�DP�҅���  ���9  �U�E؃��  ����t!�ȃ�s�M�;�w�ȃ�s�M؋}��;�v� � �U�E؍Mԃ��t�ȃ�s�M؋}��;�r�ڿ �U�E؋}�+�tz����   ����t!�ȃ�s�M�;�w�ȃ�s�M؋]��;�v蘿 �U�E؍Mԃ��t��s�E؋U��;�r�t� �EЋHLQWjV�� ��;���   �U�E؋M��AA�M�9M�u|�������}� �M�s{j j�#���������]؉]�������u��Q����u�������u��D�����uB�UЋBL�M�PQ���������t�u�M��T������'�Mԃ���E�������M��9����E��M��,�������M�d�    Y_^[�M�3�轫 ��]� �����������U���SV��F W�~@98u�}u�~< u�]K��]�~L ��   ������tw��u�}t�M�VLQSR�O� ����uX�NL�E�PQ�C� ����uD�V 9:u�N�9�V �FA�Ή�V0+ȃ�A�
�E�M��U�_�H�ND^�     �P�H[��]� �E�X{_3�^��H�H�H[��]� �������������U����EV��~L �MW�}�E��M���   ���F�����t�FL�U�RP�� ����uk��t�NLjWQ�r� ����uT�FL�U�RP�f� ����u@�M�V �ND�N@9
u�FAPPQ�������E�M��U��H�ND_�     �P�H^��]�  �E�X{_��@    �@    �@    ^��]�  �����������U��QSVW�}���    ��t�E9Fw;Fv蟼 �E�]���G9^w;^v胼 �]����t;�t�o� �G;�tB�VPRS�����؋F���E���;�t��I ���y����ǔ   ;}�u�E_�^^[��]� ��_^[��]� ����S��V�s3�;�t(W�{;�t���4����Ɣ   ;�u�CP��  ��3�_^�C�C�C[����������������SV��3�W��9^Lt�}�����u3��FLP�� ����t3��Έ^H�^A�����^L����_�^<�ND^[����U��j�hHed�    PQVW�p�3�P�E�d�    ��u��}W�L� 3�j��N��v�GR�A   �QP�U��Q������ƋM�d�    Y_^��]� �U��j�hXdd�    P��D�p�3�P�E�d�    jh(w�M��E�   �E�    �E� �Z����E�P�M��E�    �����h���M�Q�E�w詺 ��U��EVP�������w��^]� ����U��j�hHfd�    P��SVW�p�3�P�E�d�    j �M��К �=� ���E�    �]�u+j �M�譚 �=� u��@�����M�贚 �}�5��;ps"�H����u�x t�C� ;ps�P�4��3�����uN��t���F�E�WP�|��������uh<w�M��&� h��M�Q蠹 �u��Ή5���k��V覛 ���M��E������� �ƋM�d�    Y_^[��]��������������U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U��j�h�dd�    P��   SV�p�3�P�E�d�    �E3ۉ]�����   9��   j��  �����u�]���t7�M�E�P�<���P��\����E��E�   �����   �F    �$v�3��M�E�   �1��t�����\����]��]�����t�}�r�U�R�y�  ���   �M�d�    Y^[��]�U����US�]V�uW�}2��E��M��E��E�PQRWVS����+�$I�������������    +ȍ�_^[��]��������U��V�uW�};�t*S3ۃ~r�FP�߷  ���F   �^�^��;�u�[_^]����U��Q�E�V�u3҉j��N��R�A   �QP�U��Q������^��]����������U��j�h�dd�    P��SVW�p�3�P�E�d�    �e��u�}3ۉu�]���$    ;}tY�u�u��E�;�tj�S�F   �^W�Έ^�������]��u���ǋu�};�t�]V���"�����;�u�3�SS�ɶ �ƋM�d�    Y_^[��]���������������U��j�hed�    P��   �p�3�P�E�d�    �E���A�I#���   �} t	j j �\� ��t5hxw�M��s����E�P�M��E�    �@���h���M�Q�E� w�"� ��t5h`w�M��9����U�R�M��E�   ����h���E�P�E� w�� hHw��l���������l���Q�M��E�   �����h���U�R�E� w譵 �M�d�    Y��]� �����U��j�hHed�    PQVW�p�3�P�E�d�    ��u��}W�\� 3�j��N�w�GR�A   �QP�U��Q������ƋM�d�    Y_^��]� �U��EVP������� w��^]� ����U��QS3�V��WSS�^$�^�^�F  �F   �^�^�^ �.���j��  ����;�t6�� ��� j �M����(� �C���s@�C�M��<� �~$_^[��]�_�^$^[��]���������������U��j�h�fd�    PQV�p�3�P�E�d�    ��u��E�    �����P�S�  ���M�d�    Y^��]�U��j�hxed�    PQVW�p�3�P�E�d�    ��u���v�~H �E�    t�����~8�E�������u��t���f��W�ݳ  ���N蠘 �M�d�    Y_^��]��U��V���u����Et	V詳  ����^]� ���������������U��j�h�ed�    P��SVW�p�3�P�E�d�    �E�P��f��P�E�    �����}������E�������t;j �M�藓 �G��v	���sH�G�w����֍M�#�蜓 ��t
��j���Ћ�E�RP���ҋM�d�    Y_^[��]� ���U��V3�W�}��F�F�F;�u_2�^]� ��I�$	v����PW���������    +ύ��F�F_�V�^]� �����������U��j�h�ed�    P��   �p�3ŉE�SVWP�E�d�    �e��ًC��u3���K+ȸ���������������} �C  �s��+K�������ыM������º"""+Љ�p���;�s�����;��  ����"""+�;�s3���;�s��j W�?����u+s�ȸ������E������P���U������p���+ƍ�RQ���E�    �������p����E�KRPQ���d����U��p�������+ƍ��C�MRPQ���?����s�K+θ��������������E��t	V��  ����p�������+ύȋM�S����+эЉK�C�  ��p���R�ݰ  ��j j 踰 ��+M�u��������������¹   ��t����;Esy�}�E��p�������+�����QRP���~����K+M��t���P�������C��������+�WP���E�   ����s�[�E��t���R+�SP� ������N�E����+���p�����P���P+�W��������p����UQWR�C�������t���P�E�VP��������M�d�    Y_^[�M�3���� ��]� ���������������U��j�hfd�    P��<  SVW�p�3�P�E�d�    �e���u�F��u3���N+ȸ��g����������ڋ}����  �N+N���g����������¹�Ϻ+�;�s������8;��m  ���躑Ϻ+�;�s3���;�s��j S�ؿ���M+N�E츧�g����������E�i��   E�3Ƀ��M��M��MQWP���x����U�E�NRPQ���E�   �.����U�F�M�iҔ   U��E�   RPQ���	����F�N+ȸ��g�������������F�E�������t�NQP��������VR�9�  ���E�i۔   i��   ���^�~�F�M�d�    Y_^[��]� �]����u�}�~�M��i��   �PW�t�����~ �M�i��   �M�iҔ   �R�V�P���W躭  ��j j 蕭 �N+M���g�����������;���   �MQ��L���辻���E�N��i۔   �RQP���E�   ������N+M��L���R���g�����������+��FWP���E������^�v�U��L���Q+�VR�E�   �*�������L����   �E�M�i��   �Q�R�U�P�o���j j 转 �EP����������i��   �^S��+�SP���E�   �E�6����M�USQR�F����������P�E�WP�������������E������}����M�d�    Y_^[��]� ���������U��Q�M�U�E� �E�P�EQ�MR�UPQR���������]�����U��j�hHfd�    P��SVW�p�3�P�E�d�    j �M��P� �=� ���E�    �]�u+j �M��-� �=� u��@�����M��4� �}�5��;ps"�H����u�x t�Ì ;ps�P�4��3�����uN��t���F�E�WP���������uh<w�M�覧 h��M�Q� � �u��Ή5��y]��V�&� ���M��E�����蛋 �ƋM�d�    Y_^[��]��������������U��V�uW�};�tS�]j�j S���Q�����;�u�[_^]������U��Q�E�MV�uPQV�E�    ���������^��]����������U��j�h�fd�    P��SVW�p�3�P�E�d�    �e��u�}3ۉu�]���$    ;�vZ�u�u��E�;�t�Ej�S�F   �^P�Έ^����O���]��u�ǋu�};�t�]V���2�����;�u�3�SS�٩ �M�d�    Y_^[��]�U��j�h�fd�    PQV�p�3�P�E�d�    ��j�ӥ  3Ƀ�;�t�0�3���N�N�N�ƋM�d�    Y^��]��������U��j�h�fd�    PQV�p�3�P�E�d�    �M��A��P�D
��w�q����E�    ������F��H�D1�`u�M�d�    Y^��]�������������U��EVWP�����������B�����Є�t�G<    _^]� �ωw<跶��_^]� �U���   �p�3ŉE�SV�ًCW�   �u�}��{�u��+ȸ��������������;�vH9{v�T� �K+K�E�P���������������+�VWP�������_^[�M�3��A� ��]�| s]9{v�
� �K���t����M�;Kv�� �M���M�V��|�����|����������t����M���|���WPQR��t���P��������M�_^3�[�ϔ ��]�| �������������U��j�hgd�    P��SVW�p�3�P�E�d�    ��^�F�}��+ȸ��g������������E�    ;�v79^v�8� �N+N�EP���g�����������+�WSP�������PsN9^v��� �F��U�E;Fv�� �E�W�U܉M�R�M�E�������M�P� SQRP�M�Q��������M�E����������M�d�    Y_^[��] �U��E�UP��Q�MQR������]� �U��j�h8gd�    PSVW�p�3�P�E�d�    ��3�9^L��   �E�M�UPQR��� ����;���   ���FH�^A�"����O�N0�N4�G�M�F�F�~ �~$�~L��Q�ΉFD�^<豳��P�]����������B�����Є�t!�M�^<�X���ƋM�d�    Y_^[��]� �Ή~<諳���M�X���ƋM�d�    Y_^[��]� 3��M�d�    Y_^[��]� �������U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U��j�hygd�    P��4�p�3ŉE�SVWP�E�d�    �e��u�}3ۉủu��E�   �]�]ԉ]��E�;}te�uĉu��E�;�tj�S�E��F   �^P�Έ^�b���W���E��v������ũ�뻋uȋ}�;�t�]V���������;�u�3�SS荤 �}�r�M�Q藤  ���ƋM�d�    Y_^[�M�3��v� ��]�������V�qX�������V�Xu�ш ��^�����V���HW�13��@u�@(��ȋB0�Ѓ��u�   ��I΅�t�Aǃy( u��j P�E���_��^�U��QV��F��t�M�Q�N�VRQP������VR�ף  ���P�F    �F    �F    跣  ��^��]����������������U��VW�y��wX������V�Xu��� ���Et	W�s�  ����_^]� ��������U��j�h�gd�    P��SVW�p�3�P�E�d�    �e���u��H�D1΅��(  �I,��t������} ��   ��P�L2����   �MQ����XV��P�E�    �;������M���U����B�L0(�A �8 �E�   t�Q0�: ~� � ���P�҃��u!��H�D1΃��y( u��j P������W���JHu*�E�������H΃y ue��M�d�    Y_^[��]� ��H�L1(����딋M��B��H���x( u�����H�Hu�E�������>Ëu��j j �ܡ �A���y( u��j P����2��M�d�    Y_^[��]� ��������U��SVW�}���    ��t�E9Fw;Fv�p� �E�]���G9^w;^v�T� �]����t;�t�@� �O;�t5�F�E �UR�UR�URQPS������V�؋EP�NQRS�3�����(�^��_^[]� ����U��Q�UV�uW�}�E� �E�P�ER��QPVW�i�������    +΍�_^��]� ��U��SV�uW�}��+ϸ�$I�����������    +ȋE�ɋ�+�;�t+ƉE��E��V�0�/���;�u�_^��[]�����U��j�h�gd�    PQV�p�3�P�E�d�    ��u��E���Q�D(��t�H�"� �E�P�E�    ������F�ƋM�d�    Y^��]� ����U���SV��FW�E�9Fv�̟ �~�;~v轟 �M��QSWP�U�R������_^[��]������������U��j�h'hd�    P��SVW�p�3�P�E�d�    ���}�3��E�9Et��w�GXhu�E��E�   ��Q�`u�G��p����5����_j �Ή^(�F,    �����~( �F0u�F����j P���c����F    ��Q���E�   ��w�»������v�CH �CA �ͬ��3��CL���C<�KD�ǋM�d�    Y_^[��]� ������U��j�hwhd�    P��SVW�p�3�P�E�d�    ���}�3��E�9Et��w�GPhu�E��E�   ��Q�`u�G��p����5����_j �Ή^(�F,    �����~( �F0u�F����j P���c����F    ��Q�E�M��PQ���E�   ��v������ǋM�d�    Y_^[��]� �U��j�h�hd�    P��SVW�p�3�P�E�d�    �e���u�   S3�V�M��}�~�����}� �}���   �}��~{��H�L1(�A �8 �]�t�Q0�: ~� � ���P�҃��u	]��@�M;�u.^��H�L1(�Q �: t�A0�8 ~	��I ���B���
+���s�M��E�    �}�M� �~ u����J��΅�tA�y( u��j P�����E���Q�D(�E�������t�H要 �ƋM�d�    Y_^[��]� ^�M�ˉM��Q�L2(�W����'����M��@��H���x( u�����H�Hu�E�    �oDËu��?���j j �'� ����������������U��j�h�hd�    P��SVW�p�3�P�E�d�    �e��u3�WV�M܉}��E� �o����}� �}���   ��I�E�P��BO��P�E��(������M���E� �N���Mj�W�|�����B�0�A�E���~�����r������I(�A �8 t�Q0�: ~� � ���P�҅�v	���uy�M��E�    �}��@ƀ}� �@    u����I΅�t�Aǃy( u��j P�]����E܋�J�D(�E�������t�H�� �ƋM�d�    Y_^[��]ËS���JH�{����MPj������H�L1(�E�O茺���K����M��B��H���x( u�����H�Hu�E�    �:FËu�&���j j �\� �����U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U��Q�M�U�E� �E�P�EQ�MR�UPQR�;�������]�����U��QVW�}��;��W  �G�O+ȸ�$I����������Eu�������_��^��]� �NS�^+˸�$I�����������9MwY�GSP�GP�M����MQ�N�VRQP�����O+O��$I�������������    +ЋF[��_�N��^��]� ��u3���V+ӉU���$I���U��������9Ew+�G��    +э�SQP�M�����F�O�U��PQR�M��t�FPS���.����FP��  ���O+O��$I�����������P���������t�N�W�GQRP�������F[_��^��]� ������������U��j�hid�    P��X�p�3ŉE�SVWP�E�d�    �e��E��E��F�u���u�E���N+ȸ�$I����������E��}����  �^��+N��$I����������¹I�$	+�;�s������M��;��  ����I�$	+�;�s�E�    �M��ʉM�;�s�E���j Q������]+^�ȸ�$I��������3���ڋU����E��E�R��    �M�+Í�WQ�Ή]��W����U��E�NRPQ���E�   ������E�ߍ�    +Ӎ��V�EQRP���E�   ������^�N+˸�$I��������������t�VRS���H����FP���  ���E���    +ȋE�����    +ωV���V�F�  �]����u��}�~��    +ƍ�Q�M�W�������~(�U���    +ȍ���    +ƍ�RQ�M������W�z�  ��j j �U� +]��$I�����������;���   �M�Q�M�������E�N��    +��ۍRQP���E�   �����N+M�U�R��$I�����������+��FWP���E������^�v�U�M�Q+�VR�E�   ��������M��   �M��    +��M��Q���R�U�P�����j j 耕 �E�P�M������F��    +��P���P+�W���E�   �E�������M��UQWR�F�����E�P�E�SP�T������M�艿���M�d�    Y_^[�M�3��� ��]� �����������U��j�hKid�    PQV�p�3�P�E�d�    ��u��E��F�@   �@    �@ ��E�    ��t0PQ������Q���D��t�    �M�d�    Y^��]� �ƋM�d�    Y^��]� ������������U���SV��^W�~��+ϸ�$I�����������u3��3;�v�� �M���t;�t��� �M+ϸ�$I������������M�U�EQjRP���j����^;^v�ē �6W�M��u��]�������E�M��U�_^��P[��]� �����U���SVW���G��u3���O+ȸ�$I�����������_��+O��$I�����������;�s.�U�E� �M�Q�MR�GPQjS����������__^[��]� 9_v�� �U�RSP�E�P������_^[��]� ���������������U��j�h�id�    PW�p�3�P�E�d�    �}�E�E�   ;E,tP��u詒 �ML�EP�����E��u葒 �E��t#�MQP�y�����J���Dt3��E��E;E,u��}(�UL�r�EP�w�  ���}H�E(   �E$    �E r�M4Q�S�  ���ǋM�d�    Y_��]���������������U��j�h�id�    P��V�p�3�P�E�d�    �ML�UL�E� �E�P�ELQRP�� �̍U,�e�RQ�E�   �������čM�e�QP�E������u��V�E�������T�}(r�UR襑  ���}H�E(   �E$    �E r�E4P聑  ���ƋM�d�    Y^��]�������������U�����t]��]���������������̡����   ��ǀ�   `O�p   �������������������������������U��E�� t��t3�]ù�b2 �����]ø   ]����j j j jdjdhZ� j���  � ����U��j�h.jd�    PQV�p�3�P�E�d�    j j h8jH��  ���E��E�    ��t	���   �3�Pj�E������Q' ��P���H�Q`����e�V�ҡ��H�Qdj j�h`yV�҃�j j�E�   �' ��PhZ� �E������7 ��$�M�d�    Y^��]�������4 �����������U��j�h�id�    PQV�p�3�P�E�d�    ��u��R4 �N�E�    �@y�����ƋM�d�    Y^��]������������U��j�h�id�    PQV�p�3�P�E�d�    ��u��N�E�    �8������E�������3 �M�d�    Y^��]�����������U��V�������Et	V���  ����^]� ��%p�%p�%p�%p������U��E��� ]�̡����   ���   �� Q��Y�������̡��H�Qj��҃���������������U����H�U�AR�Ѓ�]��������U����H�A]����������������̡�V��H���   j�V�҃���^����U����UV��H���   RV�Ѓ���^]� �����������U���V��H���   j�V�ҡ��H�U���   j VR�Ѓ���^]� �����̡��P�BQ��Y�U����UV��H���   j VR�Ѓ���^]� ���������U����P�EP�EPQ���   �у�]� �������������U����P�EP�EP�EPQ���   �у�]� ���������U���VW���H�Qj��ҋ�����u_^]� �U���H���   RVW�Ѓ�_��^]� ����������U����P�EPQ�J�у�]� ����U����P�EPQ�J�у����@]� ��������������̡��P�BQ��Yá��P�BQ�Ѓ����������������U����P�EPQ�J�у�]� ����U����P�EPQ�Jh�у�]� ����U����P�EPQ�Jt�у�]� ����U����P�EPQ�Jl�у�]� ����U����P�EPQ�Jp�у�]� ����U����UV��H�AlRV�Ѓ����u3�^]� ���QP�B|V�Ѓ�^]� �U����P�EPQ�J|�у�]� ����U���VW�}��H�QlWV�҃����u	�E_^]� ���H�QHWV�҃�_^]� ��������������U���VW�}��H�QlWV�҃����u	�E_^]� ���H�QLWV�҃�_^]� ��������������U���VW�}��H�QlWV�҃����u�E�U_^]� ���H���   WV�҃�_^]� ��������U���VW�}��H�QlWV�҃����tI���H���   WV�ҋ�����   �QV�҃���u�����   �Q`jV�҃�_^]� �E_^]� �������������U���VW�}��H�QlWV�҃����u	�E_^]� ���H�QDWV�҃�_^]� ��������������U�����VW�}��H�QlWV�҃����u�M��E��Q�I_�P�H^��]� ���B�P`W�M�VQ�ҋ�M��P�@���Q_�A��^��]� ����������U�����0VW�}��H�QlWV�҃����u�E�u�   ���_^��]� ���H�AdW�U�VR�Ћ��E���   ���_^��]� ���������U�����VW�}��H�QlWV�҃����u0���H�u�Q`V�ҡ��H�U�ApVR�Ѓ�_��^��]� ���Q�BPWV�Ћ��Q�J`���E�P�у���t$���B�Pp�M�QV�ҡ��H�QV�҃����H�u�Q`V�ҡ��H�Ap�U�VR�Ћ��Q�Jl�E�P�у�_��^��]� �����������U�����VW�}��H�QlWV�҃����u�E�uP���b  _��^��]� ���Q�BTWV�Ѓ��M�E�fa  �E��t	P�M���c  �MQ��d  �u���U�R���a  �M���a  _��^��]� ����������U����P�EVWPQ�J\�ы��u�����B���   j�V�х�t ���B���   j VW�у�_��^]� ��_��^]� ��������������U����P�EPQ�J\�у�]� ����U�����VW�}��H�QlWV�҃����u�M��E�I_��H^��]� ���B�PXW�M�VQ�ҋ�M�@��_�A���^��]� ������U����P�EP�EPQ�J$�у�]� U����P�EP�EPQ�J(�у�]� U����P�EP�EP�EPQ���   �у�]� ���������U����E�P�EQ�$PQ�J �у�]� �������������U����E���E�   �E��B���   �U�R�URQ�Ћ����   �
�E�P�у���]� ������U����P�EP�EPQ�J<�у�]� U����P�EP�EPQ�J@�у�]� U����P�EP�EPQ�J,�у�]� U����P�EP�EPQ�J0�у�]� U����P�EP�EPQ�J8�у�]� U����P�EP�EPQ�J4�у�]� U����P�EPQ���   �у�]� �U����P�EP�EPQ���   �у�]� �������������U����P�EP�EP�EPQ���   �у�]� ���������U����P�EP�EPQ���   �у�]� �������������U����P�EPQ���   �у�]� �U����P�EPQ���   �ы����   �QXP�҃�]� ���������������U����P�EPQ���   �ыU�M��RQ���6- ]� ��U����P�EP�EP�EPQ���   �у�]� ���������U����P�EP�EPQ���   �у�]� �������������U����P�Eh#  P�EPQ���   �у�]� ��������U����P�EhF  P�EPQ���   �у�]� ��������U����P�EPQ���   �ы����   �URP�A`�Ѓ�]� �����������U����P�EPQ���   �у�]� �U����P�EP�EPQ���   �у�]� �������������U����P�EP�EPQ���   �у�]� ������������̡��P���   Q��Y��������������U��M��U�������Dz"�A�B������Dz�A�B������Dz3�]ø   ]��U����W�E��������u�   �3����U����Az�   �3�3���;���V������Au���]���E��r�$�rr �]���E����E��������z���]���E��r�$�>r ���_��^u�E������+ ��_]� ��������������U���V�u�W�}�������Dz�F�G������D{R�G����]�E�$��q �]�E�F��]�E�$�]��q �]���E�E�������D{_�   ^��]�_3�^��]�������������U���VW�M������E�}��t-���Q4P�B�Ѓ��M��u�����_3�^��]Ë�R(����H0�QW�҃��M��tԋ�R Q�MQ���ҍM���	������t���H0���   �U�RW�Ѓ��M�����_��^��]�������������U��VW�}�������=NIVb��   ��   =TCAbgtF=$'  t*=MicM��   j hIicM��������WP�B����_^]� ��BW����_�   ^]� j hdiem��������WP�B����_^]� =INIb��   �~ uŋ�B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� 聥  _3�^]� =cnys����_3�^]� ������V����y���H0�Vh�`�҉F���F    ��^�����V��F��y��t���Q0P�B�Ѓ��F    ^�����̡��P0�A���   P�у����������U����P0�E�I���   PQ�҃�]� �������������̡��I�P0���   Q�Ѓ���������̡��P0�A���   j j j j j j j j j4P�у�(������̡��P0�A���   j j j j j j j j j;P�у�(�������U����P0�E�IPQ���   �у�]� ��������������U����E V��P�M������MQh8kds�M��������E     �B0���   �M Q�M�U�R�Uj Q�MR�UQ�MR�VQj2R�Ћu ��(�M�������^��]� ������̡��I�P0���   Q�Ѓ����������U��V��F��u^]� ���Q0�M ���   j j j j j Q�Mj QjP�ҡ��H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uË��Q0P�B�Ѓ������̋A��u� ���Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5��v0Q�MQP���   R�U�R�Ћu�    �F    �����   j P�BV�Ћ����   �
�E�P�у�$��^��]� �������U����P0�E�I�R PQ�҃�]� �U��A��t)���Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�Vl�҃�^]� ����������U��y u3�]� V�u�W�}�؉��ډ���P4�A�JlWVP�ы�ډ����ى_^]� �����U��A��u]� ���Q4�M�RlQ�MQP�҃�]� ����U��A��u]� ���Q4�M�RtQ�MQP�҃�]� ����U��y u3�]� V�u�W�}�؉��ډ���P4�A�JtWVP�ы�ډ����ى_^]� �����U���VW��htniv�M������EPhulav�M������hgnlfhtmrf�M�������MQhinim�M������URhixam�M������EPhpets�M������MQhsirt�M������E �}$=  �u�����tPh2nim�M��_���Wh2xam�M��Q����E�U�RP�M�Q������������   �Q8P�ҋ�����   ��U�R�Ѓ��M��<���_��^��]�  ��U���V��htlfv�M������EQ�$hulav�M��&����EPhtmrf�M�������EQ�$hinim�M������EQ�$hixam�M�������EQ�$hpets�M�������M,Qhsirt�M��x��������E ��������Dzn���]$����Dzd�؋U(Rhdauq�M��G����M�E�PQ�U�R������������   P�B8�Ћ����   �
���E�P�у��M��1�����^��]�( ��Q�$h2nim�M��5����E$Q�$h2xam�M��!����t���������������U����S�]V�EW�}$Wj ���T$���$haerf�E ���\$�E�\$�E�\$��$P�x�������   ��MWj ���T$�$haerf�E ���\$�E�\$�E�\$�C�$Q���3�����tM��UWj ���T$���$haerf�E ���\$�E�\$�E�\$�C�$R�������t_^�   []�  _^3�[]�  ���������U���V��hCITb�M��z����EPhCITb�M������MQhsirt�M������URhulav�M������M�E�PQ�U�R�����������   P�B8�Ћ����   �
���E�P�у��M��q�����^��]� ��������U��E��Vj ��P�M�Q�M�P  �UPR���9�������H�Al�U�R�Ѓ���^��]� ����������U��E��UPj ���T$�$htemf�E���\$�E�\$�E�\$�E�$R����]� �����������U��E��Pj ���T$�U�$hrgdf�E���xy���py�����]�E�\$�E�����]�E�\$�M���]�E�\$�E�$R�%���]� �U��E��Pj ���T$�U�$htcpf�E����u�����]�E�\$�E���]�E�\$�}�]�E�\$�E�$R�����]� �������������U��Q��u3�]� �E�E�H� V�5��v0Q�MQ�M���\$�E�$QPR�V4�҃�^]� ������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�V8�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�V8�҃�^]� ����������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�V<�҃�^]� ����������U��SVW���W��t$�E�H�5��^0� �uQVP�C<R�Ѓ���u	_^3�[]� �W��t��E�H� ���[0Q�NQPR�S<�҃���t̋W��tŋE�H� �=��0Q��VP�G<R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5��v0Q�MQ�MQPR�VH�҃�^]� ������U��QV3�W��u3��,�E�H� �5��v0Q�MQPR�V8��3Ƀ�9M������U�MVR�E�����_^]� �������������U��AV��u3��"�M�Q�	�5��v0R�URQP�F8�Ѓ����M�UQ�MR������^]� ��������U��AV��u3��"�M�Q�	�5��v0R�URQP�F<�Ѓ����EQ�M�$Q�M������^]� �����U�����V���U��V�U��]�W��t$�E�H� �=��0Q�M�QPR�W<�҃���u
_3�^��]� �V��t�E�H� �=��0Q�M�QPR�W<�҃���tˋV��tċE�H� �5��v0Q�M�QPR�V<�҃���t��M�E�PQ�M�����_�   ^��]� ���U�����A�U�V�U�W�]��u3��&�M�Q�	�5��v0R�UR�U�RQP�FH�Ѓ����E�}���t�M�QP���e����E���t�EQ�$P�������_��^��]� ����U��E$�UVP�E��M Q�Mj R�UPQ�Mj R�6���P�EP���:���^]�  �����U��E,�E(�UVj P���\$���E$�M �$Q�E�M���\$�E�\$�E�\$���$R������EQ�$P�������^]�( ���U����EVQ�$��MP������]��Mj j ���T$�$htemf�E���\$�E�\$�E�\$�E�$Q���w���^]� ��U���E�EVj ���\$���E�M�\$�E�\$���$P�O���Q�M�$Q������^]� �����������U���E�EVj ���\$���E�M�\$�E�\$���$P�����Q�M�$Q�������^]� �����������U�����V�U�j �U����]���E$�M�\$�E��E �U��\$�E�$PQ�MR������M�UP�EPQR������^��]�  ����U����� V��H�A`�U�R�ЋM�E��j Q�U�RP�M�Q�M�����UPR���]�������H�Al�U�R�Ћ��Q�Jl�E�P�у���^��]� ������������U���HV��M���F  P�EP�M�Q�M����j j �U�R���?H  P�EP����������Q�Jl���E�P�у��M��DG  �M��<G  ��^��]� ���U�����EV�]���W�}����tQ�$P���h����]���M�U��E��U�P�]�Q�U�R�������N��u
_3�^��]� �U�E�r��=��0V�uV���\$�E��$P�G4RQ�Ѓ�_^��]� �������������U��E��S�م�u���H���   �҅�u[��]� VW���<y  ��htlfv�M�u�Z����E�}���]��M�]�E�$��\ �]�E�]��G�$��\ �]���E�M��}��]�E�$hulav����hmrffhtmrf�M��3����}����M�]�E�$�\ �]�E�]�G�$�\ �]���E�M��}�]�E�$hinim�4����}����M�]�E�$�K\ �]�E�]�G�$�7\ �]�E�}�]�E���$hixam�M��������Q�$hpets�M������j hdauq�M��s���Vhspff�M��e����E Phsirt�M��T����U�M�QR�E�P������������   P�B8�Ћ����   �
���E�P�у��M��>���_��^[��]� ���U��E��V���u���H���   �҅�u^��]� ���^w  �E�F��u3��"�M�Q�	�5��v0R�U�RQP�F<�Ѓ����E����y�M������]�E�\$�M��]�E�$� �����M��@�A��^��]� ����������U����E ��U�]���Vj �]�P��MQ�MR�E�PQ�M�U�R�����MP�EPQ���+���^��]� ����U�����UV�]���E�P�]��ERP������U�M�Q�MR���<�����^��]� ���U��A��u]� �M�Q�	V�5��v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� ���Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� ���Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U����P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� ���Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj=P�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5��v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M���	 �MQ�U�R�M��
 ��tm�}��E��tN�����   P�BH�ЋM��I����tQ�W�7���[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M��	 ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5��v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� ���Q0�M�RTQ�MQ�MQP�҃�]� U��A��u]� ���Q0�M�RXQ�MQ�MQ�MQ�MQ�MQP�҃�]� ���̋A��uË��Q0P�Bh�Ѓ�������U��A��u]� ���Q0�M�R\Q�MQP�҃�]� ����U��A��u]� ���Q0�M�R`��   �QP�҃�]� ��U��A��u]� ���Q0�M�R`QP�҃�]� ��������U��A��u]� ���Q0�M�RdQ�MQ�MQ�MQP�҃�]� ������������U���V�u�VW���H4�R�ЋE�F    �~�H� ���R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� ���Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I���R0P�EPQ���   �у�]� ������̡��I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u�� ���R0�I�RPV�uVP�EPQ�҃�^]� �����������U����P0�E�I�RtP�EP�EP�EP�EPQ�҃�]� �U����P0�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U��E�P� V�5��v0R�UR�UR�UR�URP�A�NxP�у�^]� ��������U��E� ���R0j j j j j j j P�A���   jP�у�(]� �����������U��E� ���R0j j j j j jj P�A���   jP�у�(]� �����������U��E� ���R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M������E�H� ���R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R������M��������^��]� ����������U��E�P� V�5��v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5��v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5��v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5��v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U����P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U����UVj j j j j R��H0�E�Vj P���   jR�Ћ��Q0�E�N���   PQ�҃�0^]� ���������������U����P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡��P0�A���   j j j j j j j j jP�у�(�������U����P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡��P0�A���   j j j j j j j j j(P�у�(�������U����P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U����P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡��P0�A���   j j j j j j j j jP�у�(������̡��P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}�M���tj j��������u��tj j�����������H0�U��B�IpVWP�у�_^[��]� ���������U����P0�E�I���   P�EP�EPQ�҃�]� �����̡��P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V����y���H0�Vh�`�҉F3��F�F����y�F   ��^�������V��F��y��t���Q0P�B�Ѓ��F    ^������U��E�UVj P�E��MQRPj j ���]�����t�~ t
�   ^]� 3�^]� ��U��E�A�I��u3�]� ���B0Q�H�у�]� ����U��S�]V�������=ckhc��   tu=cksatY=TCAb��   Wj hdiem�����������PSW���F   �҃~ ��t��t��u3�������P�[���_^��[]� �~ tK��B����^[]� �~ t6���������t+�F    ^�   []� =atnit�MQS������^[]� ^3�[]� ���������U��V��~ ��   W�}����   �$����E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN���M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W�|  ���F    _^]� ��Ѝލ�����,�����U��V��~ �"  �EW�}�E����   �$�����E������A��   �   ���E��������   �   ���E��������   �v���E������A��   �b�E������A��uP��������   �E�E��������u3������A{}�,�E���������E������A�����E������DzU����ء��U�H0�F���   j j j j j j j RjP���E�U��(R���\$�E�$W�9{  ���F    _^]� �ڎ���0�M�f�r�~�����U���E�E�Uj���\$�E�\$�E�$PR�w���]� ���U���E�E�Uj���\$�E�\$�E�$PR�G���]� ���U���E�E�Uj���\$�E�\$�E�$PR����]� ��̋�3�� �y�H�H�H�������������VW��3���y9~u���H4�V�R�Ѓ��~�~_^����U����P4�E�I�RxPQ�҃�]� �U��U��t3�A���I0R���   P�ҋ��Q0�M���   QP�҃�]� ���P0�E�I���   PQ�҃�]� ���̡��P4�A�JP�у������������̡��P4�A�JP�у������������̡��P4�A�JP�у������������̡��P4�A���   P�у���������̡��P4�A���   P�у����������U����P4�E�I�RP�EP�EP�EPQ�҃�]� �����U����P4�E�I�RP�EP�EP�EPQ�҃�]� �����U����P4�E�I�R PQ�҃�]� �U����P4�E�I�R$PQ�҃�]� �U����P0�E�I���   P�EP�EP�EPQ�҃�]� ��U����P4�E�I���   PQ�҃�]� ��������������U����P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U����P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U����P4�E�I�R(PQ�҃�]� �U����P4�E�I�R,P�EP�EPQ�҃�]� ���������U����P4�E�I�R0P�EPQ�҃�]� ������������̡��P4�A�J4P��Y��������������U���S�]VW3���~Pj�ˉE�E��}���j j�ˉE��o����E���H0�UR�W�E�P�ApR�Ћ��Q4�F�JP�ы��J0j �U�R�U�R�U�R�U�RP�F�P�AxR�Ѓ�,�} _^[t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ���������U����P4�E�I�R8PQ�҃�]� �U����P4�E�I�R<PQ�҃�]� �U����P4�E�I���   P�EPQ�҃�]� ���������̡��P4�A�J@P�у�������������U����P4�E�I�RDP�EPQ�҃�]� �������������U����P4�E�I�RHP�EPQ�҃�]� �������������U����P4�E�I�RLP�EPQ�҃�]� �������������U����P4�E�I�RPP�EPQ�҃�]� �������������U���VW�}��H�QW�҃���t���H4�U�ER�VP�ATWR�Ѓ�_^]� ��������������U����P4�E,P�E(P�E$P�E �IP�E�RXP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U����P4�E�I�R\P�EP�EP�EPQ�҃�]� ����̡��P4�A�JdP��Y�������������̡��P4�A�JhP�у�������������U����P4�E�I�R`P�EP�EP�EP�EP�EPQ�҃�]� �������������U����P4�E�I�RlP�EPQ�҃�]� �������������U��V�uW��t��؉�}��t��ډ���P4�A�JlWVP�у���t��ډ��t��ى_^]� �U��V�uW��t��؉�}��t��ډ���P4�A�JtWVP�у���t��ډ��t��ى_^]� �U����P4�E�I�RtP�EPQ�҃�]� �������������U���$V��~ ��   ���V�H4�AR�Ѓ} t#���Q0���   P�F�HQ�҃�^��]� ��hARDb�M܉E��E�    �y���P�M�Q�N�U�R�8��������   ��U�R�Ѓ��M�躹��^��]� ���U����P4�E�I�RpPQ�҃��   ]� ������������U����E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U����P4�E�I���   P�EP�EPQ�҃�]� �����̡��P4�A���   P�у���������̸   ����������̸   �����������U���V��H4�V�A$h�  R�Ћ��Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U����P4�E�I�R|P�EP�EP�EPQ�҃�]� �����U����P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}�M���tj j���Q�����u��tj j���=�������H4�U��B�ItVWP�у�_^[��]� ���������U��QSVW�}���3�苸��=INIb�   ��   =SACbwt+=$'  t
=MicM�Q  ��P$W����_�   ^��[��]� 3��E��E��@�MQ�U�R���Ѕ�t���E�Q4�M�P�FQ�JP�у�_�   ^��[��]� =ARDb��   j j���V���j j�ϋ��I���j j�ωE��;���j j�ωE�-����M���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>������P���h���P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� j hIicM���d����WP�B ����_^[��]� U����P4�E�I�RXh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M�躴�����Q4�JpP�FP�у��M�����^��]��������V����y���H0�Vh�`�҉F���F    �z�F   ��^��������V��F��y��t���Q0P�B�Ѓ��F    ^������U��VW�}����ϵ��=cksat`=ckhct�EPW�������_^]� �Fj j j j j j �F   ���Q0���   j j j P�у�(��t'_�F    �   ^]� �~ t��B����_^]� _3�^]� �����������U����H��H  ]��������������U����H0���   ]��������������U����H0�U�E��VWRP���   �U�R�Ћ��Q�u���B`V�Ћ��Q�BpVW�Ћ��Q�Jl�E�P�у�_��^��]������������U����H0���   ]��������������U����H0���   ]��������������U��Ej0P�"f  ��]��������������U��Ej0P��  ��P��e  ��]�����U��E�M��j0PQ�U�R��  ��P��e  ���H�Al�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P��  ��P�e  ���Q�Jl�E�P�у���]��U��Ej$P�be  3Ƀ�������]����U��Ej$P���  ��P�9e  3Ƀ�������]�����������U��E�M��Vj$PQ�U�R��  ��P��d  ��3Ƀ��B�Pl����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P���  ��P�d  ��3Ƀ��B�Pl����M�Q�҃���^��]����U����H�U�E��  RPj �у�]���������������U����H�U�ER�UP��  Rj �Ѓ�]�����������U����P4�E�I�R,P�EP�EPQ�҃�]� ���������U����P4�E�I�R0P�EPQ�҃�]� ������������̡��P4�A�J4P��Y��������������U���VW�}j ��j������j j�ωE��
����E���H0�UR�V�E�P�ApR�Ћ��Q0�E�H� �RxQ�M�Q�M�Q�M�Q�M�Q�NPQ�҃�(�} _^t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ���U��ESVW�؅�u�Y�}j hdiuM���=�������t3;3u	_^3�[]� j hIicM������;�uj h1icM��課���uӉ3_^�   []� ��������U���V�uhfnic���:�����tj
���ݰ�����uShfnic�E�P��訵���uP��������M��������.������t���"�����uhfnic���2����MQj
��蕷��^��]�U����P0�E�IP�EP�EP�EPQ���   �у�]� ��U����P0�E�IV�p� ���   V�uj j j V�uVj Pj>Q�҃�(^]� ����U����P0�E�IV�p� ���   V�uV�uj j j�Vj Pj>Q�҃�(^]� ���̡��I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V����y���H0�WVh�`�ҋ}���F�Ej hmyal���F    �F   �4z�F�@����F��t��t�F    j hhfed�������F_��^]� ���U��VW�}���菮��=ytsdt�EPW������_^]� ���Q0�F���   P�ы�B������_�   ^]� ����������3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ���������������������U��E3�h�����h  ���P�Ej BR�Uj PR�����]� �U��S�]$V�EW�}�S�]j ����T$���$�E htemf���\$�E�\$�E�\$�E�$P�r�������   �G�M�]S��j ���T$�$�E htemf���\$�E�\$�E�\$�E�$Q���'�����t:�E �US���\$���E�\$�E�\$�G�$R������t_^�   []�  _^3�[]�  U���E �ES�]VW�}$W���\$���E�\$�E�\$��$P������th�E �MW���\$�E�\$�E�\$�C�$Q���������t:�E �UW���\$���E�\$�E�\$�C�$R������t_^�   []�  _^3�[]�  ������U���E �ES�]VW�}$W���\$���E�\$�E�\$��$P�������th�E �MW���\$�E�\$�E�\$�C�$Q��������t:�E �UW���\$���E�\$�E�\$�C�$R������t_^�   []�  _^3�[]�  ������U��Q��u3�]� �E�H� V�5�W�}Q�MQ�}�v0PR�VD�ҋ�����tD�E��t=���QWP�Bp�ЋE����t#���Q��P�Bl�Ћ��Q�BW�Ѓ�_��^]� ������U�����V��H�A`�U�R�ЋU���M�QR���D�������u���H�Al�U�R�Ѓ�3�^��]� �M�Q�M�u  ���B�Pl�M�Q�҃���^��]� �������U�����V��H�A`�U�R�ЋU���M�QR��������M���E�PQ�M�B������B�Pl�M�Q�҃���^��]� ����U���V��M���  �M�E�PQ��� ����M�U���ERP�����M��  ��^��]� �������������U��EVj ��MP�L����Mh���h  �j j jj PQ��莼��^]� ���������U�����V�U�j �U����]���E$�M�\$�E��E �U��\$�E�$PQ�MR蟫���M�UP�EPQR���k���^��]�  ����U�����V�U�j �U����]���E$�M�\$�E��E �U��\$�E�$PQ�MR�?����M�UP�EPQR�������^��]�  ����U�����V�U�j �U����]���E$�M�\$�E��E �U��\$�E�$PQ�MR�ߪ���M�UP�EPQR���;���^��]�  ����U���4���H�Q`SVW�}W�ҋu��3�SS�Ή]�"���Sj�ΉE�������;��   �} ~d���H�A`�U�R�Ћ��Q�Jdj j��E�h�zP�ы��B�HW�ы��J�U�RP�A0W�Ћ��Q�Jl�E�P�у�(���B0�M����   VQ�U�R�Ћ��Q�J`���E�P�ы��B�Pp�M�QV�ҡ��H�Al�U�R�Ћ��Q�BW�Ћ��Q�R0�M�QPW�ҡ��H�Al�U�R�Ћu�E��0j ��
S������j �KQ�ΉE�����������������_^[��]���U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj AQj R�UR��譹��^]� ��������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR�o���^]� ����������U��E�E$3҃8��R�U(R�U���\$�E �$R�E���\$�E�\$�E�\$�@�E�$P����]�$ ��������������U��E�@3҃8�]��E��Rj ���T$�$htemf�E���\$�E�\$�E�\$�E�$P豹��]� �������������U��E�E3҃8��R���\$�E�\$�E�\$�@�E�$P�ڼ��]� ������U��E�E3҃8��R���\$�E�\$�E�\$�@�E�$P�
���]� ������U��E3҃8��R�UR�UR�UR�UP�EPR����]� U��E�E 3҃8��R�U���\$�E�\$�E�$P�EP�ERP�����]� �U��E�E 3҃8��R�U���\$�E�\$�E�$P�EP�ERP����]� �U��E�E 3҃8��R�U���\$�E�\$�E�$P�EP�ERP�U���]� �U��E�E 3҃8��R�U���\$�E�\$�E�$P�EP�ERP�����]� �U��E3҃8V�u��V��RP�EP�����^]� ����������U��Q��u3�]� �E�E�H� V�5��v0Q�MQ�M���\$���E�$QPR�V4�҃�^]� ���U��EVj ��MP���������u�    �F^]� ��u9Ft�   ^]� ���U��EVj ��MP��������u�    �F^]� ��u9Ft�   ^]� ���U����EVQ�$��MP�����]����u�E�    �^^]� ��u�F�E������D{�   ^]� ���������������U���$��VW�U����U��M�]�E�PQ�M�U�R�Ǥ����x��@�U�}�E����u�V�~_�    �F^��]� ��u�E�P�NQ藬������t�   _^��]� ��U�����V���]��M��E��]�PQ�M�U�R�Y������@�U��E���u�    �V�F^��]� ��u�E�P�NQ�#�������t�   ^��]� ���������������U���VW�}�M�;}u\�uj htsem���\�����uGPhrdem���K�����u6�E�E��EP�M�Q�M�}��޹����t�U�M�R�.  _�   ^��]� _3�^��]� �������U���VW�}�M�;}u\�uj htsem���ܡ����uGPhrdem���ˡ����u6�E�E��EP�M�Q�M�}�讹����t�U�M�R�  _�   ^��]� _3�^��]� �������U���SVW�}��;}ua�uj htsem���\�����uLPhrdem���K�����u;��E��E�]P�M�Q�M�}��l�����t�EQ���$�Z  _^�   [��]� _^3�[��]� �U���(�ESW�}�M�;�t;Et	;E��   �]j htsem���̠������   Phrdem��跠����uv�E��M�U��U��U�R�]؉E�M�E�P�M�Q�M�U�R�E�    �E�    �}��E�    ������t+�M؋U܃��ĉ�M��P�H�M���  �   _[��]� _3�[��]� ���U���SVW�}��;}uk�uj htsem��������uVPhrdem���������uE��M�E��]���E�P�]�Q�M�U�R�}��������t�E��M�PQ���  _^�   [��]� _^3�[��]� �������U�����0VW���H�A`�U�R�Ћ��Q�J`�E�P�ыE���U�RP�M�Q�M輡�����J�U�RP�Ap�Ћ��Q�Jl�E�P�ы��B�Pl�M�Q�ҡ��H�Q`��V�ҡ��H�Ap�U�VR�Ѓ����  ���Q�Jl�E�P�у�_^��]� ������������U���SVW�}��;}ul�uj htsem��謞����uWPhrdem��蛞����uF���H�A`�U�R�Ѓ��M�Q�M�U�R�}��E�    ������U��u���H�AlR�Ѓ�3�_^[��]� ����R�j�����T  ���H�Al�U�R�Ѓ�_^�   [��]� ��U��V�u����  ��^]� �����������U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�A�E������D{�   ]� ���������U��V�����u�E�M�U�F�N�    �V^]� ��u�EP�NQ�Ŧ������t�   ^]� ���U��V�����u�E�M�    �F�N^]� ��u�UR�FP�{�������t�   ^]� ���������U��V��F��y��t���Q0P�B�Ѓ��E�F    t	V�'  ����^]� ��������������U��V��~ ��yu���H4�V�R�Ѓ��E�F    �F    t	V�A'  ����^]� �������U���V��3ɍF��H��������M��M����   �RQ�M�QP�ҡ����   ��U�R�Ѓ���^��]��������������U��V�����u �    ���H�Ap���UVR�Ѓ��(��u$���Q�R P�EP�NQ�҃���t�   ���H�Al�UR�Ѓ�^]� ��U����P�EP�EP�EPQ�Jd�у�]� �����������̡��H$�Q�����U����H$�U�AR�Ѓ�]��������U����H$�A]����������������̡�V��H$�QDV�҃���^���������U���V��H$�QDV�ҡ��U�H$�AdRV�Ѓ���^]� U���V��H$�QDV�ҡ��U�H$�ARV�Ѓ���^]� U���V��H$�QDV�ҡ��H$�U�ALVR�Ѓ���^]� ���P$�BHQ��Y�U����P$�EPQ�JL�у�]� ���̡��P$�BQ�Ѓ����������������U����P$�EP�EP�EPQ�J�у�]� ������������U����P$�EP�EP�EPQ�J�у�]� �����������̡��P$�BQ�Ѓ����������������U���VW�}��H�Q`W�ҡ��H$�QV�ҋ�����t ���H�QpWV�ҡ��H�QV�҃���_^]� ���������U����P$�EPQ�J�у�]� ���̡��P$�B(Q��Yá��P$�BhQ��Y�U����P$�EPQ�J,�у�]� ����U����P$�EPQ�J0�у�]� ����U����P$�EPQ�J4�у�]� ����U����P$�EPQ�J8�у�]� ����U����UV��H$�ALVR�Ѓ���^]� ��������������U����H$�QDV�uV�ҡ��H$�U�ALVR�Ћ��E�Q$�J@PV�у���^]���������������U����UV��H$�A@RV�Ѓ���^]� ��������������U����P$�EPQ�J<�у�]� ����U����P$�EPQ�J<�у����@]� ���������������U��V�u���t���Q$P�B�Ѓ��    ^]���������U����P$�EP�EPQ�JP�у�]� U����P$�EPQ�JT�у�]� ���̡��H$�QX�����U����H$�A\]�����������������U����P$�EP�EP�EPQ�J`�у�]� �����������̡��H(�������U����H(�AV�u�R�Ѓ��    ^]��������������U����P(�EP�EP�EP�EP�EP�EPQ�J�у�]� ���P(�BQ�Ѓ����������������U����P(�EPQ�J�у�]� ����U����P(�EP�EP�EPQ�J�у�]� ������������U����P(�EP�EPQ�J�у�]� U����P(�EjP�EPQ�J�у�]� ��������������U����P(�EP�EPQ�J�у�]� ���P(�B Q�Ѓ���������������̡��P(�B$Q�Ѓ���������������̡��P(�B(Q�Ѓ����������������U����P(�EPQ�J,�у�]� ����U����P(�EPQ�JP�у�]� ����U����P(�EPQ�JT�у�]� ����U����P(�EPQ�JX�у�]� ����U����P(�EPQ�J\�у�]� ����U����P(�EPQ�J`�у�]� ����U����P(�EPQ�Jp�у�]� ����U����P(�EPQ�Jd�у�]� ����U����P(�EPQ�Jh�у�]� ����U����P(�EPQ�Jl�у�]� ����U�����V���E�    �E�    �H(�A`�U�RV�Ѓ�����   �E���uI���Q�J`�E�P�ы��B�M�@pQ�U�R�Ћ��Q�Jl�E�P�у��   ^��]� ���J��H  j j P�҃��E���u���H(�Q,j�V�҃�3�^��]� ���Q(�M��Rj QPV�҃���u�E�P��  ��3�^��]� �M��U�j IQ�MR�����E�P��  ���   ^��]� ���U�����V��H�A`�U�R�Ѓ��M�Q������^��u���B�Pl�M�Q�҃�3���]� ���H$�E�I�U�RP�ы��B�Pl�M�Q�҃��   ��]� �U��Q���P(�E�PQ�JP�у���u��]� �E3�8U���   ��]� �����U���VW�}��H(�QhWV�҃���t$���H(�Qh��WV�҃���t_�   ^]� _3�^]� ����U���VW�}��H(�QhWV�҃���t>���H(�Ah�WRV�Ѓ���t%���Q(�Bh��WV�Ѓ���t_�   ^]� _3�^]� ����������U���VW�}��H(�QlWV�҃���t>���H(�Al�WRV�Ѓ���t%���Q(�Bl��WV�Ѓ���t_�   ^]� _3�^]� ����������U��VW�}W��������t8�GP��������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U����P(�EPQ�J0�у�]� ����U����P(�EPQ�J4�у�]� ����U����P(�EPQ�J8�у�]� ����U����P(�EPQ�J<�у�]� ����U����P(�EPQ�J@�у�]� ����U����P(�EP�EPQ�Jt�у�]� U����P(�EPQ�JD�у�]� ����U����E�P(�BHQ�$Q�Ѓ�]� �U����E�P(�BL���$Q�Ѓ�]� ��������������̡��H,�Q����̡��P,�B8�����U����H,�A V�u�R�Ѓ��    ^]�������������̡��P,�B<�����U����P,�R@��VW�E�P�ҋu�����H$�QDV�ҡ��H$�QLVW�ҡ��H$�AH�U�R�Ѓ�_��^��]� �������U����P,�E�RH��VWP�E�P�ҋu�����H�Q`V�ҡ��H�QpVW�ҡ��H�Al�U�R�Ѓ�_��^��]� ��̡��H,�j j �҃��������������U����P,�EP�EPQ�J�у�]� U����H,�AV�u�R�Ѓ��    ^]�������������̡��P,�BQ�Ѓ���������������̡��P,�BQ�Ѓ���������������̡��P,�BQ�Ѓ���������������̡��P,�B,����̡��P,�BD����̡��P,�B0�����U����P,�R4]�����������������U����H,�A$]�����������������U����H,�AL]�����������������U����H,�A(]�����������������U���VW�}��H$�QDW�ҡ��H,�QV�ҋ�����t ���H$�QLWV�ҡ��H$�QV�҃���_^]� ���������U����H�I]�����������������U����H�A]�����������������U����H�I]�����������������U����H�A]�����������������U����H�I]�����������������U����H��\  ]��������������U����H�A ]�����������������U����H�A$]�����������������U����H�I,]�����������������U����H��p  ]��������������U����H��t  ]��������������U����H��x  ]��������������U����H$�QDVW�}W�ҡ��H�Q(���ҋ���t ���H$�QLWV�ҡ��H$�QV�҃���_^]���������������U����H$�QDVW�}W�ҡ��H��X  ���ҋ���t ���H$�QLWV�ҡ��H$�QV�҃���_^]������������U����H��d  ]��������������U����H�U��L  ��VWR�E�P�ы��u���B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�҃�_��^��]����������������U��V�ujV��������^]���������̡��H���   ��U����H���   V�uV�҃��    ^]�������������U����P�EP�EP�EPQ���   �у�]� ��������̡��P���   Q�Ѓ������������̡��P���   Q�Ѓ�������������U����P�EPQ�JL�у�]� ����U����P�EPQ�JP�у�]� ����U����P�EPQ�JT�у�]� ����U����P�EPQ�JX�у�]� ����U����P�EPQ�J\�у�]� ����U����P�EPQ�J`�у�]� ����U����P�EPQ���   �у�]� �U����P�EPQ�Jd�у�]� ����U����P�EPQ�Jh�у�]� ����U����P�EPQ�Jl�у�]� ����U����P�EPQ�Jp�у�]� ����U����P�EPQ�Jt�у�]� ����U����P�EPQ�Jx�у�]� ����U����P�EPQ�J|�у�]� ����U����P�EPQ���   �у�]� �U����P�EPQ���   �у�]� �U����P�EPQ���   �у�]� �U����P�EPQ���   �у�]� �U����P�EP�EPQ���   �у�]� �������������U����P�EP�EPQ���   �у�]� �������������U����P�EPQ���   �у�]� �U��E��t ���R P�B(Q�Ѓ���t	�   ]� 3�]� U����P �E�RhQ�MPQ�҃�]� U��E��u]� ���R P�B,Q�Ѓ��   ]� ������U����P�EPQ�
�у�]� �����U����P�EPQ�J�у�]� ����U����P�EPQ�J�у�]� ����U����P�EPQ�J�у�]� ����U����P�EPQ�J�у�]� ����U����P�EPQ�J�у�]� ����U����P�EP�EPQ���   �у�]� �������������U����E�P�BQ�$Q�Ѓ�]� �U����E�P�B���$Q�Ѓ�]� ���������������U����P�EPQ�J �у�]� ����U����P�EPQ�J$�у�]� ����U����P�EPQ�J(�у�]� ����U����P�EPQ�J,�у�]� ����U����P�EPQ�J0�у�]� ����U����P�EPQ�J4�у�]� ����U����P�EPQ�J8�у�]� ����U����P�EPQ�J<�у�]� ����U����P�EP�EP�EP�EPQ���   �у�]� �����U����P�EPQ�JD�у�]� ����U����P�EPQ���   �у�]� �U����P�EP�EPQ�JH�у�]� ���P���   Q�Ѓ�������������U����P�EPQ���   �у�]� �U����P�EPQ���   �у�]� �U����P�EPQ���   �у�]� �U����P�EP�EPQ���   �у�]� ������������̡��P���   Q�Ѓ�������������U����P�EP�EPQ���   �у�]� ������������̡��P���   Q�Ѓ������������̡��P���   Q�Ѓ������������̡��P���   Q�Ѓ�������������U����H���   ]��������������U����H���   ]��������������U����H�U�E��VWRP��4  �U�R�Ћ��Q�u���B`V�Ћ��Q�BpVW�Ћ��Q�Jl�E�P�у�_��^��]������������U����H��8  ]��������������U���VW�}��H$�QDW�ҡ��H$�Q V�ҋ�����t ���H$�QLWV�ҡ��H$�QV�҃���_^]� ���������U���VW�}��H$�QDW�ҡ��H$�Q$V�ҋ�����t ���H$�QLWV�ҡ��H$�QV�҃���_^]� ���������U���V�uV�E�P�������e������Q$�JH�E�P�у���^��]� �������U����P(�} ����PQ�J0�у�]� �������������U���VW�}���H(�]�E�QHQ�$V�҃���t-�G���H(�]�E�QHQ�$V�҃���t_�   ^]� _3�^]� U���VW�}���H(�]�E�QHQ�$V�҃���tO�G���H(�]�E�QHQ�$V�҃���t-�G���H(�]�E�QHQ�$V�҃���t_�   ^]� _3�^]� ��������������U���VW�}���H(�QL���$V�҃���tG���G�H(�QL���$V�҃���t)���G�H(�QL���$V�҃���t_�   ^]� _3�^]� ����������U��VW�}W���������t8�GP���������t)�OQ���������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W��������t8�GP��������t)�O0Q���������t��HW���������t_�   ^]� _3�^]� ������������U���S�]VW���H�QPj S�ҋ���H��H  j Fj V�҃��E��u���H(�Q,j�W�҃�_^3�[]� ���Qj VP�BTS�Ћ��Q(�B@VW�Ѓ���t"���E�Q(�JVPW�у���t�   �3��UR��  ��_��^[]� ����U���V�E���MP����P���#������Q�Jl���E�P�у���^��]� ���U���V�u�E�P���������Q$�J�E�P�у���u���B$�PH�M�Q�҃�3�^��]á��H�A�U�jR�Ѓ���u�M�Q��������t����H�QjV�҃���u0���H�Q V�҃���u���H$�AH�U�R�Ѓ�3�^��]Ë��Q$�JH�E�P�у��   ^��]�������U���<� SVW�E�    ��t�E�P�   ����������Q$�JD�E�P�   �у��u����B$�}�HDW�ы��B$�HLWV�у���t���B$�PH�M�Q����҃���t���H$�AH�U�R�Ѓ���_^[��]����U��V�u���t���QP�B�Ѓ��    ^]���������U����H��  ]��������������U��E��t�x��u�   ]�3�]������U��E��s�   VW�xW� ������u_^]Ã} tWj V��  ��_������F��   ^]����������������U����E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�| ������u_^]�Wj V�&�  ��_������F��   ^]�������������U����E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�� ������u_^]�Wj V��  ��_������F��   ^]�������������U����E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�| ������u_^]�Wj V�&�  ��_������F��   ^]�������������U����E��t#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   VW�xW�� ������u_^]�Wj V��  ��_������F��   ^]���������U�����tO�} �Et#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËM�UQR�7�����]���U����E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW� ������u_^]�Wj V��  ��_������F��   ^]�������������U����E��t#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   VW�xW� ������u_^]�Wj V�2�  ��_������F��   ^]���������U�����tO�} �Et#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËM�UQR�������]���U��M��t.�=� t�y���A�uP�  ��]á��P�BQ�Ѓ�]�������U��M��t.�=� t�y���A�uP���  ��]á��P�BQ�Ѓ�]�������U��M��t.�=� t�y���A�uP��  ��]á��P�BQ�Ѓ�]�������U��M��t.�=� t�y���A�uP�Q�  ��]á��P�BQ�Ѓ�]�������U��M��t.�=� t�y���A�uP��  ��]á��P�BQ�Ѓ�]�������U��M��t.�=� t�y���A�uP���  ��]á��P�BQ�Ѓ�]�������U��M��t.�=� t�y���A�uP��  ��]á��P�BQ�Ѓ�]�������U��M��t.�=� t�y���A�uP�Q�  ��]á��P�BQ�Ѓ�]�������U����H|�]����H|�h   �҃�������������U��V�u���t���Q|P�B�Ѓ��    ^]���������U����P|�EP�EPQ�J�у�]� U����P|�EP�EPQ�J�у�]� U����P|�EP�EPQ�J�у�]� U����P|�EPQ�J�у�]� ���̡��HL��8  ��U����H@�AHV�u�R�Ѓ��    ^]�������������̡��HL�������U����H@�AHV�u�R�Ѓ��    ^]�������������̡��PL���   Q�Ѓ�������������U����PL�EP�EPQ���   �у�]� �������������U���V��HL���   V�҃���u���U�HL���   j RV�Ѓ�^]� �����   �ȋBP�Ћ����   �MP�BH��^]� �����̡��PL��p  Q�Ѓ�������������U����PL�EP�EPQ��t  �у�]� ������������̡��HL�Q�����U����H@�AHV�u�R�Ѓ��    ^]��������������U��V�uW������l�����U�HL�AVRW�Ѓ�_��^]� �U����PL�EPQ��   �у�]� �U����PL�EP�EPQ�J�у�]� ���PL�B Q�Ѓ���������������̡��PL�B$Q�Ѓ���������������̡��PL�B(Q�Ѓ����������������U����PL�EP�EPQ�J,�у�]� U����PL�EPQ��|  �у�]� �U����PL�EP�EP�EPQ�J0�у�]� ������������U����PL�EP�EP�EP�EPQ�J4�у�]� �������̡��PL�B8Q�Ѓ���������������̡��PL�B<Q�Ѓ����������������U����PL�EP�EPQ��`  �у�]� ������������̡��PL���   Q�Ѓ�������������U����PL��VQ��   �E�P�ыu��P���6k���M��nk����^��]� �����U����PL�E��T  ��VPQ�M�Q�ҋu��P����j���M��*k����^��]� ̡��PL�B@Q�Ѓ���������������̡��PL�BDj Q�Ѓ��������������U����PL���   ]��������������U����PL���   ]��������������U����PL��4  ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL��  ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL��0  ]��������������U����PL�EPQ�JT�у�]� ���̡��PL�BQ��Y�U����PL�EP�EPQ�JX�у�]� U����PL�Ej PQ�J\�у�]� ��U����PL�Ej PQ�J`�у�]� ��U����PL�EjPQ�J\�у�]� ��U����PL�EjPQ�J`�у�]� ��U���SVW3��E��P�M��}��}��E��  �}�}��A  W�M�Q�U�R����G  ���M�����3  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U���3�V�E�E�E��P�M��E�   �E�   �E��  �^@  j�M�Q�U�R���MG  �M��3  �����   ��U�R�Ѓ�^��]�����������U������UVW3���}��}����   �I(R�E�P�у��U�R�M��E��  �}�}���?  j�E�P�M�Q����F  �M��2  �����   ��M�Q�҃�_^��]� ��U������UVW3���}��}����   �I(R�E�P�у��U�R�M��E��  �}�}��Z?  j�E�P�M�Q���IF  �M��2  �����   ��M�Q�҃�_^��]� ��U���SVW3��E��P�M��}��}��E��  �}�}���>  W�M�Q�U�R����E  ���M����1  ��t+�u���I��������   ��U�R�Ѓ�_��^[��]� �����   �JL�E�P�ыu��P�����������   ��M�Q�҃�_��^[��]� ���U���SVW3��E��P�M��}��}��E��  �}�}��4>  W�M�Q�U�R���E  ���M�����0  ��t+�u�����������   ��U�R�Ѓ�_��^[��]� �����   �JL�E�P�ыu��P������������   ��M�Q�҃�_��^[��]� ���U���SVW3��E��P�M��}��}��E��  �}�}��t=  W�M�Q�U�R���DD  ���M����'0  _^��[t�����   ��U�R�������]Ë����   �J<�E�P���]������   ��M�Q���E�����]���������������U���SVW3��E��P�M��}��}��E��  �}�}���<  W�M�Q�U�R���C  ���M����w/  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U���SVW3��E��P�M��}��}��E��  �}�}��<  W�M�Q�U�R����B  ���M�����.  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�@�u������   �
�F�E�P�у�_��^[��]� �̡��PL��  Q��Y��������������U����PL�E��  ��jPQ�M�Q�ҋ�M�@�A�������]� �������U����PL�E��  ��j PQ�M�Q�ҋ�M�@�A�������]� �������U���SVW3��E��P�M��}��}��E��  �}�}��:  W�M�Q�U�R���A  ���M����g-  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�@�u������   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}���9  W�M�Q�U�R����@  ���M����,  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�@�u������   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��49  W�M�Q�U�R���@  ���M�����+  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�@�u������   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��t8  W�M�Q�U�R���D?  ���M����'+  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U����E3�V�]��E�E�E��P�M��E�   �E��  �7  j�M�Q�U�R���>  �M��v*  �����   ��U�R�Ѓ�^��]� ���������U����EV��M�E�3�Q�M��E�   �E��  �E�E��O7  j�U�R�E�P���>>  �M��*  �����   �
�E�P�у�^��]� ��������U������UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}���6  j�E�P�M�Q���=  �M��)  �����   ��M�Q�҃�_^��]� ��U������UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��J6  j�E�P�M�Q���9=  �M��)  �����   ��M�Q�҃�_^��]� ��U������UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}���5  j�E�P�M�Q���<  �M��(  �����   ��M�Q�҃�_^��]� ��U������UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��J5  j�E�P�M�Q���9<  �M��(  �����   ��M�Q�҃�_^��]� ��U����EV��M�E�3�Q�M��E�   �E��  �E�E���4  j�U�R�E�P����;  �M��'  �����   �
�E�P�у�^��]� ��������U���SVW3��E��P�M��}��}��E��  �}�}��t4  W�M�Q�U�R���D;  ���M����''  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�@�u������   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��3  W�M�Q�U�R���:  ���M����g&  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U���SVW3��E��P�M��}��}��E��  �}�}��3  W�M�Q�U�R����9  ���M����%  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U������UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��2  j�E�P�M�Q���	9  �M���$  �����   ��M�Q�҃�_^��]� ��U����EV��M�E�3�Q�M��E�   �E��  �E�E��1  j�U�R�E�P���8  �M��f$  �����   �
�E�P�у�^��]� ��������U����EV��M�E�3�Q�M��E�   �E��  �E�E��?1  j�U�R�E�P���.8  �M���#  �����   �
�E�P�у�^��]� ��������U����H���   ]��������������U����H���   ]�������������̡��H���   ����H���   ��U����H���   V�u�R�Ѓ��    ^]�����������U����H���   ]��������������U����HL�QV�ҋ���u^]á��H�U�ER�UP��@  RV�Ѓ���u���Q@�BHV�Ѓ�3���^]����������U����H�U�E��@  R�U�� P�ERP�у�]������U����H���   ]��������������U����H�U0�E,R�U(P�E$R�U P�ER�Uj P�ER�UP�ER�UP���   R�Ѓ�0]����������̡��PL�BdQ�Ѓ���������������̡��PL�BhQ�Ѓ����������������U����PL�EP�EPQ�Jl�у�]� U����PL�EPQ��d  �у�]� �U����PL�EPQ��  �у�]� ̡��PL�BtQ�Ѓ����������������U����PL�EP�EP�EPQ���   �у�]� ���������U����PL�EP�EP�EPQ�J|�у�]� ������������U���<��SV��HL�QW�ҋ�3ۉ}�;��w  �M��!U���M�E�Qh]  �ȉ]ȉ]Љ]ԉ]؉]��E�   �]��}ĉE��/]�������   �PSSW���҅���   ���HL�Q W�ҋ���;���   ��    �����   �B(���ЍM�Qh�   ���u��  ������   �M�;���   �����   ���   S��;�tm�����   �ȋB<V�Ћ����   ���   �E�P�у�;�t���B@�HHV�у���;��]����}��M��S���M��T����_^[��]� �}����B@�HHW�ы����   ���   �M�Q�҃��M��:S���M��BT��_^3�[��]� ������̡��PL���   Q�Ѓ������������̡��PL���   Q�Ѓ�������������U����PL�EPQ���   �у�]� ̡��PL���   Q�Ѓ�������������U����PL�EPQ���   �у�]� �U����PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U�E�EVh��h��h��h��R�Q�UR�UR�UQ�A�$�5��vLRP���   Q�Ѓ�,^]� ������������̡��PL���   Q�Ѓ�������������U����PL�EPQ���   �у�]� �U����PL�EPQ���   �у�]� �U����PL�EPQ���   �у�]� �U����PL�EPQ���   �у�]� �U����PL�EPQ���   �у�]� ̡��PL��<  Q�Ѓ�������������U����PL�EP�EP�EPQ��h  �у�]� ���������U����PL�EP�EP�EP�EP�EPQ��@  �у�]� �U����PL�EP�EP�EPQ��D  �у�]� ���������U����PL�EP�EP�EP�EPQ��H  �у�]� �����U����HL��$  ]��������������U����HL��(  ]��������������U����HL��,  ]�������������̡��HL��\  ��U���(��V3��u؉u܉u��u�u�u�u��E�   �u􋈜   ���   W�ҋ}�E�;�t`;�t\���QLjP���   ���ЋM��U�Rh=���M�}��  �������   ���   �U�R�Ѓ��M؉u���N����_^��]Ë����   ���   �E�P�у��M؉u��N��_�   ^��]����������U���(��V3��u؉u܉u��u�u�u�u��E�   �u􋈜   ���   W�ҋ}�E�;�t`;�t\���QLjP���   ���ЋM��U�Rh<���M�}��9  �������   ���   �U�R�Ѓ��M؉u��N����_^��]Ë����   ���   �E�P�у��M؉u���M��_�   ^��]���������̡��H8�������U����H8�AV�u�R�Ѓ��    ^]��������������U����P8�EP�EPQ�J�у�]� U����P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U����P8�EP�EPQ�J�у�]� U����P8�EP�EP�EP�EP�EPQ�J�у�]� ����U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H�A0]�����������������U����H�I4]�����������������U����H�Q`V�uV�ҡ��H�Q<V�҃���^]�����̡��H�Q@�����U����H�ID]����������������̡��H�QH����̡��H�QL�����U����H�AP]�����������������U����H�AT]�����������������U����H���  ]��������������U����H��|  ]��������������U����H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡��H���   ����H��   ��U����H�U�ER�UP�ER�UP���   Rh�*  �Ѓ�]����������������U����H�A]�����������������U����H�Ad]�����������������U����H�Ah]�����������������U����H�Al]����������������̡��H�Qp����̡��H�Qt����̡��H�Qx�����U����H�A|]�����������������U����H���   ]��������������U����H���   ]��������������U����H���  ]��������������U����H��X  ]��������������U����H���   ]��������������U����H���  ]��������������U��V�u��袱�����H�U���   VR�Ѓ���^]������U����H���   ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]�������������̡��H���   ��U����H���  ]��������������U����H��P  ]��������������U����H��T  ]��������������U��V�u���"H�����H���   V�҃���^]���������̡��H���  ��U����H��\  ]��������������U����H�U���   ��R�E�P�ы�M��P�@�Q�A������]�������U����H��  ]��������������U��U�E���H�E���   R���\$�E�$P�у�]�U����H���   ]��������������U����H��   ]��������������U����H��h  ]��������������U����H��l  ]��������������U����H��  ]��������������U����H���  ]��������������U����H��$  ]��������������U����H��(  ]��������������U����H��,  ]��������������U����H��0  ]��������������U����H��4  ]��������������U����H��8  ]��������������U����H��<  ]��������������U����H��@  ]��������������U����P���E�P�E�P�E�PQ��D  �у����#E���]����������������U����P���E�P�E�P�E�PQ��D  �у����#E���]����������������U����P���E�P�E�P�E�PQ��D  �у����#E���]����������������U����H���  ]��������������U��V�u(V�u$�E�@���R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@���R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U����P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U����P0�EP�EP�EP�EPQ���   �у�]� ����̡��P0���   Q�Ѓ�������������U����P0�EP�EPQ���   �у�]� �������������U����P0�EP�EP�EP�EPQ���   �у�]� ����̡��P0���   Q�Ѓ������������̡��H0���   ��U����H0���   V�u�R�Ѓ��    ^]�����������U����H���  ]��������������U����H���  ]�������������̡��H���  ����H��  ��U����H��,  ]��������������U����H��8  ]��������������U����H��0  ]��������������U����H��(  ]��������������U����H��H  ]��������������U����H�U�E���  ��VR�UPR�E�P�ыu�    �F    �����   �Qj PV�ҡ����   ��U�R�Ѓ� ��^��]��������U���Vj hLGOg�M��JA��P�E�hicMCP�k������M��A�������   �JT�E�P�у���u(�u����@�������   ��M�Q�҃���^��]á����   �AT�U�R�Ћu��P����@�������   �
�E�P�у���^��]�������������U����H��`  ]��������������U����H���  ]��������������U����H�U���  ��V�uVR�E�P�у��������M�������^��]�����U����H���  ]��������������U����H�U���  ��VWR�E�P�ы��u���B�H`V�ы��B�HpVW�ы��B�Pl�M�Q�҃�_��^��]����������������U����H�U���  ��VWR�E�P�ы��u���B�H`V�ы��B�HpVW�ы��B�Pl�M�Q�҃�_��^��]����������������U����H���  ]��������������U����H���  ]��������������U����H��   ]��������������U����H��  ]��������������U����H��  ]��������������U��E�M�U��VWPQR�����     �@    �����   �M�Rj QP�ҡ��H���  �U���R�Ћ��Q�u���B`V�Ћ��Q�BpVW�Ћ��Q�Jl�E�P�у�(_��^��]�����������U����H�U�E��  ��VR�UPR�E�P�ыu�    �F    �����   �Qj PV�ҡ����   ��U�R�Ѓ� ��^��]��������U���  �p�3ŉE��M�EPQ������R��  ���H���  ������Rh�z�ЋM�3̓��<�  ��]�������������U����H��h  ��V�U�WR�Ћ��Q�u���B`V�Ћ��Q�BpVW�Ћ��Q�Jl�E�P�у�_��^��]����U����H��l  ��V�U�WR�Ћ��Q�u���B`V�Ћ��Q�BpVW�Ћ��Q�Jl�E�P�у�_��^��]����U����H���  ���҅�tbh���M��)<���EPh���M��XD���MQh���M��GD��j �U�R�E�hicMCP�#��������   �
�E�P�у��M��D<����]�U����H���  ��V�҅�u���H�u�Q`V�҃���^��]�Wh!���M��;���EPh!���M��C��j �M�Q�U�hicMCR���������   P�BH�Ћ��Q�u���B`V�Ћ��Q�BpVW�Ћ����   �
�E�P�у�$�M��;��_��^��]�����������U����H���  ���҅�u��]�Vh#���M���:���EPh#���M��C��j �M�Q�U�hicMCR����������   P�B8�Ћ����   �
���E�P�у��M���:����^��]������U����H���  ���҅�u��]�Vhs���M��D:���EPhs���M��sB��j �M�Q�U�hicMCR�O��������   P�B8�Ћ����   �
���E�P�у��M��\:����^��]������U����H��,  ]��������������U����H���  ]��������������U����H��0  ]��������������U��V�u���t���QP���  �Ѓ��    ^]������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]�������������̡��H���  ��U����H���  ]��������������U����H���  ]�������������̡��H���  ��U����H�U���  ��VR�E�P�ыu��P���38���M��k8����^��]�����U����H���  ]��������������U����H��   ]��������������U����H��  ]��������������U����H��  ]��������������U����H��  ]��������������U����H��  ]��������������U���h����M��7��j �E�P�M�hicMCQ�9��������   ��M�Q�҃��M��Z7����]�������U����H��   ]��������������U����H���  ]��������������U����H��L  ]�������������̡��H��P  ��U����H��T  ]������������������������������U����H��|  ]��������������U����H�A`�U��� R�Ћ��Q�Jdj j��E�h�zP�ыUR�E�P�M�Q�mt�����B�Pl�M�Q�ҡ��H�A�U�R�Ћ��Q�Jl�E�P�у�,��]��h�PhD ��q  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h�jhD ��p  ����t
�@��t]��3�]��������Vh�j\hD ����p  ����t�@\��tV�Ѓ���^�����Vh�j`hD ���p  ����t�@`��tV�Ѓ�^�������U��Vh�jdhD ���ip  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�jhhD ���)p  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh�jlhD ����o  ����t�@l��tV�Ѓ�^�������U��Vh�h�   hD ���o  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h�   hD ���fo  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�jphD ���o  ����t�@p��t�MQV�Ѓ�^]� � ^]� ��U��Vh�jxhD ����n  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�jxhD ���n  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�jxhD ���Yn  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� ������������̋���������������h�jhD ��m  ����t	�@��t��3��������������U��V�u�> t+h�jhD ��m  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h�jhD �m  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�jhD ���9m  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�jhD ����l  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�j hD ���l  ����t�@ ��tV�Ѓ�^�3�^���Vh�j$hD ���l  ����t�@$��tV�Ѓ�^�3�^���U��Vh�j(hD ���Yl  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�j,hD ���	l  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�j(hD ����k  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�j4hD ���|k  ����t�@4��tV�Ѓ�^�3�^���U��Vh�j8hD ���Ik  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�j<hD ����j  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh�jDhD ���j  ����t�@D��tV�Ѓ�^�3�^���U��Vh�jHhD ���j  ����t�M�PHQV�҃�^]� U��Vh�jLhD ���Yj  ����u^]� �M�PLQV�҃�^]� �����������U��Vh�jPhD ���j  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�jThD ����i  ����u^Ë@TV�Ѓ�^���������U��Vh�jXhD ���i  ����t�M�PXQV�҃�^]� U��Vh�h�   hD ���vi  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�h�   hD ���&i  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�h�   hD ����h  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ���h  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ���Vh  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ���h  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh�h�   hD ��g  ����u���H�u�Q`V�҃���^��]ËM���   WQ�U�R�Ћ��Q�u���B`V�Ћ��Q�BpVW�Ћ��Q�Jl�E�P�у�_��^��]��U��Vh�h�   hD ���Fg  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�h�   hD ����f  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   hD ���f  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   hD ���vf  ����t���   ��t�MQ����^]� 3�^]� �Vh�h�   hD ���9f  ����t���   ��t��^��3�^����������������U��Vh�h�   hD ����e  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�h�   hD ���e  ����t���   ��t�MQ����^]� ��������U��Vh�h�   hD ���fe  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������VW��3����$    �h�jphD �e  ����t�@p��t	VW�Ѓ��� �8 tF��_��^�������U��SW��3�V��    h�jphD �d  ����t�@p��t	WS�Ѓ��� �8 tkh�jphD �d  ����t�@p��tWS�Ѓ����� h�jphD �^d  ����t�@p��t�MWQ�Ѓ��� �;uG�c����E^��t�8��~=h�jphD �d  ����t�@p��t	WS�Ѓ��� �8 u_�   []� _3�[]� U��Vh�j\hD ����c  ����t3�@\��t,V��h�jxhD �c  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�j\hD ���ic  ����t3�@\��t,V��h�jdhD �Gc  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�j\hD ���c  ����tG�@\��t@V�ЋEh�jdhD �E��E�    �E�    ��b  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�j\hD ���b  ����t\�@\��tUV��h�jdhD �gb  ����t�@d��t
�MQV�Ѓ�h�jhhD �>b  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�j\hD ����a  ������   �@\��t~V��h�jdhD ��a  ����t�@d��t
�MQV�Ѓ�h�jhhD �a  ����t�@h��t
�URV�Ѓ�h�jhhD �a  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh�jthD ���Fa  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�j`hD �a  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh ���_�����^��]� ������U���Vh�h�   hD ���`  ����tR���   ��tH�MQ�U�R���ЋuP������h�j`hD �z`  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t�����   P�B@��]� �E��t�����   P�BD��]� �����   R�PD��]� �����U����P@���   ]��������������U����P@���   ]��������������U����P@���   ]��������������U����P@���   ]��������������U������   ���   ]�����������U������   ���   ]����������̡��P@���   ����P@���   ��U����P@���   ]�������������̡��P@���   ������   �Bt��U����P@���   ]�������������̡��P@���   ��U����P@���   ]��������������U���V��H@�Q$V�ҋM����t��#������Q@P�B V�Ѓ�^]� �̡��PH���   Q�Ѓ�������������U����P@�EPQ���   �у�]� ̡��P@���   Q�Ѓ������������̡��P@�B,Q�Ѓ����������������U����P@�EPQ�J(�у�]� ����U����P@�EP�EP�EPQ�JP�у�]� ������������U����P@�EPQ�JT�у�]� ����U����P@�EP�EPQ�JX�у�]� U����P@�EPQ�J\�у�]� ����U������   �R]��������������U������   �R]��������������U������   �R ]��������������U������   ���   ]�����������U����E���   �E���   P�EP�EQ�$P�EP�EP��]� �����������U������   ���   ]����������̡����   �B$����H@�Ql�����U����H@�Apj�URj �Ѓ�]����U����H@�Apj�URh   @�Ѓ�]�U����H@�U�E�IpRPj �у�]�̡����   ����U��V�u���t�����   P�B�Ѓ��    ^]�����̡����   �Q ��U��V�u���t�����   P�B(�Ѓ��    ^]�����̡��H@�Ql�����U��V�u���t���Q@P�BH�Ѓ��    ^]���������U����H@���   ]��������������U��V�u���t���Q@P�BH�Ѓ��    ^]��������̡��PH���   Q�Ѓ�������������U����PH�EPQ���  �у�]� �U����H �Id]�����������������U��}qF u?V�u��t6�����   �BDW�}W���ЋM���B@VQ�HhW�у����(��_^]���̡��P@���   ��U����P@���   ]��������������U����P@���   ]�������������̡��P@���   ��U��Q���P�EWP�M�Q�JP�ы�����u_��]� ���B��H  SVj �_j S�ы�����u	^[_��]� �M���B�U��@TQSVR�Ѓ��> ��^[_��]� ���������������U����H�Q`VW�}W�ҡ��H�U�ADR�Ћ�����t"���Q�BpWV�Ћ��Q�BV�Ѓ���_^]���������U����H�Q`V�uV�ҡ��H�U�E�I|VRP�у���^]��������������U����H�Q`VW�}W���E���H�U�E��R�UP�ERPQ�I@�$�ы�����t"���B�HpWV�ы��B�HV�у���_^]���U����p�3ŉE�V�uW�}�E�0�E�x�   �   ��    ��������
s0�7�D�B��y���D� �H�Q`W�ҡ��H�Adj j��U�RW�ЋM�����_3�^���  ��]�������U��� V�uW�}���&  ��   @vp���H�A`�U�R�Ћ��Q�Jdj j��E�h�zP�у��U�Rj0j jj �ǋֱ�ڹ  �U�E�m��z�]�EQ�E��$P�x�������   ����   ��   v`���H�A`�U�R�Ћ��Q�Jdj j��E�h�zP�у��U�Rj0j jj �ǋֱ
�X�  �U�E�m��z�]�E�y�����|6��   v,j h�z�M������mPj0��zj jj �]�E�?���j h�z�M������P�E�WP�
������uPV��W�����Q�Jl�E�P�ы��B�Pl�M�Q�҃�_��^��]���������������U����PT�EP�EPQ�J�у�]� U����PT�EPQ�J8�у�]� ����U����PT�EPQ�J@�у�]� ����U����PT�E�Rh��PQ�M�Q�ҋ�M��P�@�Q�A������]� ������U����HT�U�j R�Ѓ�]�������U����H@�AHV�u�R�Ѓ��    ^]�������������̡��HT�j hG  �҃�����������U����H@�AHV�u�R�Ѓ��    ^]��������������U����HT�U�j R�Ѓ�]�������U����H@�AHV�u�R�Ѓ��    ^]��������������U����E�PH�B Q�$Q�Ѓ�]� �U����PH�EPQ���   �у�]� �U����PH��0VWQ�JP�E�P�ы��E���   ���_^��]� �������������U����PH��0VWQ�JT�E�P�ы��E���   ���_^��]� �������������U����PH�EPQ���  �у�]� �U����PH�EPQ��   �у�]� �U����PH�EP�EPQ��D  �у�]� �������������U����PH�EP�EPQ��H  �у�]� ������������̡��PH���  Q�Ѓ�������������U����PH�EPQ���  �у�]� ̡��PH�Bdj Q�Ѓ��������������U����PH�EPj Q�Jh�у�]� �̡��PH�BdjQ�Ѓ��������������U����PH�EPjQ�Jh�у�]� �̡��PH�BdjQ�Ѓ�������������U����PH�EPjQ�Jh�у�]� ��U����PH�EP�EPQ���   �у�]� �������������U����PH�EP�EPQ���   �у�]� ������������̡��PH�BtQ�Ѓ����������������U����PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���p-  ������t�E���QH���   PVW�у���_^]� �����U��EVW���MPQ��-  ������t�M���BH���   QVW�҃���_^]� ̡��PH��  Q�Ѓ������������̡��PH��  Q�Ѓ�������������U����PH�EPQ��  �у�]� �U����PH�EPQ��  �у�]� �U����PH�EP�EPQ��P  �у�]� �������������U����PH�EP�EPQ��  �у�]� ������������̡��PH���  Q�Ѓ������������̡��PH���  Q�Ѓ������������̡��PH���  Q�Ѓ������������̡��PH��   Q�Ѓ������������̡��PH��$  Q�Ѓ�������������U����PH�EP�EPQ��(  �у�]� �������������U����PH�EP�EP�EPQ��,  �у�]� ���������U����PH�EPQ��<  �у�]� ̡��PH��t  Q�Ѓ�������������U����PH�EP�EPQ��@  �у�]� �������������U����PH�EPQ��h  �у�]� ̡�V��H@�QhWV�҃�j h�  ����������HH���   h�  V�҃���
��t_3�^Ë�_^��������������̡��P@�BhQ�Ѓ�j h�  ������U����E�PH�E��,  ��P�EPQ�$Q�M�Q�ҋ�M��P�@�Q�A������]� ��������U����E�PH�E��0  ��P�EPQ�$Q�M�Q�ҋ�M��P�@�Q�A������]� ��������U����PH�EP�EPQ��4  �у�]� ������������̡��PH��8  Q��Y��������������U����E�PH��<  Q�$Q�Ѓ�]� �������������̡��PH��@  Q�Ѓ�������������U����PH�EP�EPQ��D  �у�]� �������������U����E�PH�EP�EQ�$PQ��H  �у�]� �����̡��PH���  Q�Ѓ������������̡��PH��L  Q�Ѓ������������̋��     �������̡��PH����  jP�у���������U����UV��HH���  R��3Ƀ������^��]� ��̡��PH����  j P�у��������̡��PH��h  Q�Ѓ������������̡��PH��l  Q�Ѓ������������̡��PH��p  Q�Ѓ�������������U����PH��Q��t  �E�P�ы�M��P�@�Q�A������]� ������̡��PH��x  Q�Ѓ�������������U����PH�EPQ��|  �у�]� �U����E�PH���  Q�$Q�Ѓ�]� ��������������U����E�PH���  Q�$Q�Ѓ�]� ��������������U����E�PH���  Q�$Q�Ѓ�]� ��������������U����PH�EPQ���  �у�]� �U����E�HH�U�ER�UP�EQ�$R�UP���   R�Ѓ�]��������������U����E�HH�U�ER�UQ���   �$P�ERP�у�]��U���E�M��z蜕  �M;�|�M;�~��]�����������U����HH�U�ER�UP���   R�Ѓ�]������������̡��PH���   Q��Y�������������̡��PH���   Q�Ѓ������������̡��PH���   Q��Y��������������U����PH�EP�EPQ���   �у�]� �������������U����PH�EP�EP�EP�EP�EPQ���  �у�]� ̋�� �z�@    ���z���Px�A�JP��Y��������U���V��Hx�V�AR�ЋE����u
�   ^]� ���Qx�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË��QxP�B�Ѓ�������U����Px�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U����E�HH�U�ER�UQ�$P���  R�Ѓ�]������U����HH���  ]��������������U����HH���  ]��������������U����E(�HH�U,�E$R�U Q�$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�(]��������������U����HH���  ]��������������U����E�PH�EPQ�$Q���  �у�]� ����������U���SV���1  �؉]����   �} ��   ���HH���  j h�  V�҃��E��u
^��[��]� �MW3��}��P  ����   �]��I �E�P�M�Q�MW�  ��ta�u�;u�Y�I ������u�E�������L�;Ht-���Bx�S�@����QR�ЋD������t	�M�P��  F;u�~��}��MG�}��  ;��v����]�_^��[��]� ^3�[��]� ��������������U�����SV�ًHH���  j h�  S�]��ҋ�����u
^3�[��]� �E��u���HH���  �'��u���HH���  ���uš��HH���  S�ҋȃ��E��t�W��  ���HH���   h�  S3��҃����  ���_�u����    ���Hx�U�B�IWP�ы�������   ���F�J\�UP�A0R�Ѓ���t�K�Q�M�  ���F�J\�UP�A0R�Ѓ���t�K�Q�M�|  �E��;Pt&�F���Q\�J0P�EP�у���t	�MS�L  ���v�B\�M�P0VQ�҃���t�M�CP�#  ���QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U����HH��  ]�������������̡��PH��  Q��Y��������������U����HH���  ]��������������U��Q��V�uW�}Q�$V���v
���]��E��E������Au������E������{����]Q�E���$V�~��_^��]���������U��� ��V�u�U�W�U��}�]�E�PV�M�Q���W
���E��E�����E��Au���U��������z�����U����E�������z���U�����]���������Au@�����U����E�������z0�����]�U��ER�]�V�E����]��E��]��?��_^��]��]�����������Au����������U����HH�U�j R�Ѓ�]�������U����H@�AHV�u�R�Ѓ��    ^]�������������̡��HH�j h�  �҃�����������U����H@�AHV�u�R�Ѓ��    ^]��������������U����HH�Vj h  �ҋ�������   �EPh�  ��  ����t]���QHj P���   V�ЋMQh(  �  ����t3���JH���   j PV�ҡ����   �B��j j���Ћ�^]á��H@�QHV�҃�3�^]�����U����H@�AHV�u�R�Ѓ��    ^]��������������U����HH�Vj h�  �ҋ�����u^]á��HH�U�E��(  RPV�у���u���B@�HHV�у�3���^]�����U����H@�AHV�u�R�Ѓ��    ^]��������������U����HH�I]�����������������U����H@�AHV�u�R�Ѓ��    ^]��������������U����PH�EPQ���  �у�]� �U����PH�EPQ���  �у�]� ̡��PH���  Q�Ѓ�������������U����HH���  ]��������������U����E�HH�U(�E$R�U P�ER�UP�ER�U���\$�E�$P��p  R�Ѓ�$]������������̡��PH��  Q�Ѓ�������������U����PH�EP�EPQ��  �у�]� ������������̡��PH��8  Q�Ѓ�������������U����PH�EP�EP�EPQ��   �у�]� ��������̡��PH��$  Q�Ѓ������������̡��PH��(  Q�Ѓ�������������U����PH�EPQ��0  �у�]� �U����PH�EPQ��4  �у�]� ̋������������������������������̡��HH��  ��U����HH��  ]��������������U����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��  �у�0]�, ���������U����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��x  �у�0]�, ���������U����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��  �у�0]�, ���������U����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��|  �у�0]�, ��������̡��PH��X  Q�Ѓ�������������U����PH�EPQ���  �у�]� ̡��PH���  Q�Ѓ�������������U����HH��\  ]��������������U����HH��d  ]��������������U�����W���HH���   j h�  W�҃��} u�   _��]� Vh�  �?  ������tq���HH���   j VW�҃��M������EPh�  �M��6���EQ�$h�  �M�������Q@�Jdj �E�PV�у��M��R���^�   _��]� ^3�_��]� �����������U��S�]�; VW��u7���U�HH���   RW�Ѓ���u���QH���   jW�Ѓ���t�   �����   ���QH���   W�Ѓ��} u(���E�QH�M���  P�ESQ�MPQW�҃��B�u��t;���U�HH�ER�USP���  VRW�Ћ����   �B(�����Ћ���uŃ; u���QH���   W�Ѓ���t3���   �W��u1���QH���   �Ћ��E�QH���   PW�у�_^[]� ���BH���   �у��} u0���M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ���QH�j h  �Ћ؃���u_^[]� �����   �u�Bx���Ћ����   P�B|���Ѕ�t_���$    ����E�QH�MP�Ej Q���  VPW�у���t�����   �ȋBHS�Ћ����   �B(���Ћ���u�_^��[]� ��U��EV���u���HH���  �'��u���HH���  ���u���HH���  V�҃���u3�^]� P�EP������^]� ���������U���@���HH���   SV�uWh�  V�ҋ����HH�Q|3�Sh�  V�}��]��҉E�3����E�E��E�;���  �����   �B���Ћ�=�  �  �QH�Bx3�Wh:  V�Ћ��QH�E䋂�   h�  V�Ћ��QHW�؋B|h�  V�]ԉ}��Ћ��QH�E苂8  V�Ћ��QH�EЋ�$  V�Ѓ�(�E��E��z��~{�M���M܋MЅ�tMj�W��N  ���t@�@�Ẽ|� ��~����%�������;�u/���hW  ;E�~�E؋��)W  E���E܋;Pu�E���E��E�G;}�|��}� tm�}�j V���S  ����   ����  ��tM���  �]�;�uB���H��H  �<[j ��j W�҃��E����   �M�WP�  P���������]���H��H  �<[3�S��SW�҃��E�;�tr�M�;�t;�tWQP��z  ���E�;�~!���QS��SP��H  �Ѓ��E�;�t4���E��QH��(  j�PV�у���t�}�;�tAjV���\  ��u'�U�R�����E�P�����M�Q�݁����_^3�[��]Ë���  �E���]����BH�H|Sh�  V�у�3�9]ԉE�]���  �}���I �MЅ��  j�S��L  �����  �@�Ẽ|� ���U�~�
���%�������;��  3�3�9J�M���   �����������tz�]��U���������M���ʋ���]��U��҉T��]�@�U؋Q�T��]��U�@B�T��Q�]�@�T��U؋]�@���T��I�U�@�L��M؋U�@@�����U�@�M�A;J�M��e����E܅��h  �+�j��P�E�P�M��7  �M�v���E��E�3�+��E����    �}� �M����E�t-�M�@���MĉU؋U�ʋU؋��U؋R�Q�U؋R�Q;]܋U��@����M؋M���U؋R�Q�U؋R�Q}j����    �E��M�9�uU�ыL�����������w4�$��`�M����4�"�U����t��M����t�
�U����t��;]�|��E�F;]��"����S  ��M�3�;G�Å���   �E��v���W��R�����Q�P�I�H�O��I�M����P�Q���P�I�H��@�E���U��Lv�����P�Q�@�A��t&�G�U�@���U��Lv	�����P�Q�@�A�G��U��@���U�v�����P�Q�@�A�G��w��U��@���U�F�v�����P�Q�@�A��w��U�F�@���U�v�����P�Q�@�A�7F��t+�G�U��@���U�v�����P�Q�@�A�wF���O�]�C��;]ԉ]�������U�R�~���E�P�~�����  ���   �B����=  ��  ���QH�B|j h(  V�Ћ��QH�����   h(  V�ЋЃ�3��U؅�~�ǅ�t�|� t�K��\K�@;�|�]��]����Q��H  �[j ��j S�Ѓ��E�����   �}� t��t�M�SQP��u  ���]؋��B��H  �j ��j S�у��E��tP��t��tSWP�u  ���M����+��RH��PQ�E���  V�Ѓ���u�M�Q��|���U�R��|����_^3�[��]á��HH�Q|j h�  V�҉E����HH�Q|j h(  V��3�3�3ۃ�9U؉Eĉ}̉]���   �u荛    �ޅ���   ���E�    ~g�u�<�R��   ����d$ �u��>��\>��EԉY�v�q�u��\7�t7�Y�^���Y�v�]�q�u�B@B����;�|��}̃|� tO�Eԋu�8�E��I���R�4����A�F�I�N�M��u���B�R�4����A�F�I�N�u�B<މ}�C;]؉]������M�3�3�;�~�Uĉt���   @;�|�U�R�b{�����E�P�V{����_^�   [��]ÍI K\V\b\n\����U��E� �M+]� ���������������U��V��V��z���Hx�AR�Ѓ��Et	V�������^]� ����������U����H ���   ]��������������U����H@�AHV�u�R�Ѓ��    ^]�������������̡��H �������U��V�u���t���Q P�B�Ѓ��    ^]���������U����P �EPQ�JP�у�]� ����U����P �EPQ�J�у�]� ����U����P �EPQ�J�у�]� ���̡��P �BQ��Y�U��V�uW�����/������H �Q VW�҃�_��^]� �����U����P �EPQ�J$�у�]� ���̡��P �BDQ�Ѓ���������������̡��P �BLQ�Ѓ����������������V����-����z�F    ��^��������U��E�A�   ]� ��������������U��E�M� P   �P   �   ]� ��� �������������V��W�~���R-��3��G��z��F�F_��^�����������V����t���Q P�B4�Ѓ��N^�,-��������������U��E��S�]V��F�K�N��u^[��]�, W�}(�v��tj�U�R�FP�ˉ}��E�    �% ���K�]0�FS�],���R SW�}$W�} W�}W�}W�}W�}WP�FQ�J0P�у�03҅���_�^[��]�, ���U���V��> t6�M��*���hNIVb�M��������H ��I8j �U�RP�у��M�����^��]��������U����t*�y t$�y t���Q �M�R8Q�MQP�҃�]� 3�]� �������U��V��FW�}��t&���t �x t�x t���P �B8jWQ�Ѓ��MQW���6��_^]� �������U��V���+���Et	V�{������^]� ��������������̡��H\�������U����H\�AV�u�R�Ѓ��    ^]�������������̡��P\�BQ��Yá��P\�BQ�Ѓ���������������̡��P\�BQ�Ѓ����������������U����P\�EPQ�J�у�]� ����U����P\�EP�EPQ�J�у�]� U����P\�EPQ�J�у�]� ���̡��P\�B Q�Ѓ����������������U����P\�EPQ�J$�у�]� ����U����P\�EP�EPQ�J(�у�]� U����P\�EP�EP�EPQ�J,�у�]� ������������U����P\�EPQ�J4�у�]� ����U����P\�EPQ�JD�у�]� ����U����P\�EPQ�JH�у�]� ���̡��P\�B8Q�Ѓ����������������U����P\�EP�EPQ�J<�у�]� U����P\�EPQ�J@�у�]� ����U���SVW�}��j �ωu���i�����H\�QV�҃���S����i��3���~=��I ���H\�U�R�U��EP�A,VR�ЋM��Q���i���U�R���i��F;�|�_^[��]� ���������������U���VW�}�E��P���(f���}� ��   ���Q\�B V�Ѓ��M�Q���f���E���t]S3ۅ�~H�I �UR����e���E�P����e���E;E�!�����Q\P�BV�ЋE@��;E��E~�C;]�|�[_�   ^��]� _�   ^��]� ���PD�BQ�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�BPQ�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ����������������U����PX��Q�
�E�P�ы�M��P�@�Q�A������]� �����������U����PX��Q�J�E�P�ы�M��P�@�Q�A������]� ����������U����PX��Q�J�E�P�ы�M��P�@�Q�A������]� ����������U����PX��0VWQ�J�E�P�ы��E���   ���_^��]� �������������U����PX��0VWQ�J�E�P�ы��E���   ���_^��]� �������������U����PX�EPQ�J�у�]� ����U����PX�EPQ�J�у�]� ����U����PX�EPQ�J�у�]� ����U����PX�EPQ�J �у�]� ����U����PX�EPQ�J8�у�]� ����U����PX�EPQ�J(�у�]� ����U����PD�EP�EPQ�J,�у�]� U����HD�U�j j R�Ѓ�]�����U����H@�AHV�u�R�Ѓ��    ^]��������������U����HD�U�j j R�Ѓ�]�����U����H@�AHV�u�R�Ѓ��    ^]��������������U����U�HD�E�	Rj P�у�]���U����H@�AHV�u�R�Ѓ��    ^]��������������U����HD�U�j j R�Ѓ�]�����U����H@�AHV�u�R�Ѓ��    ^]��������������U��U���HD�Rj h'  �Ѓ�]��U����H@�AHV�u�R�Ѓ��    ^]�������������̡��HD�j j h�  �҃���������U����H@�AHV�u�R�Ѓ��    ^]�������������̡��HD�j j h:  �҃���������U����H@�AHV�u�R�Ѓ��    ^]��������������U���3��E��E������   �R�E�Pj�����#E���]�̡��HD�j j h�F �҃���������U����H@�AHV�u�R�Ѓ��    ^]�������������̡��HD�j j h�_ �҃���������U����H@�AHV�u�R�Ѓ��    ^]��������������U��E����u��]� �E����E�    ���   �R�E�Pj������؋�]� ̡��PD�BLQ�Ѓ����������������hPh�f ��  ���������������U���Vhh�   h�f ���  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vhh�   h�f ���&  ����t���   ��t�M�UQ�MRQ����^]� U���Vhh�   h�f ����  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vhh�   h�f ���V  ����t���   ��t�M�UQ�MRQ����^]� U��Qhh�   h�f �  ����t���   �E���t�EP�U�����]�� {��]�������������U���hh�   h�f ��  3Ƀ�;�tK9��   tC�E���   ���M��$Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]ËE�   � �  �P�P�H�H�H��]��U��hh�   h�f �9  ����t���   ��t]��]����U��hh�   h�f �	  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��hh�   h�f �  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��hh�   h�f �I  ����t���   ��t]�����]�U���Vhh�   h�f �  ����tZ���   ��tP�M�UWQR�M�Q�Ћ��u���B�H`V�ы��B�HpVW�ы��B�Pl�M�Q�҃�_��^��]á��H�u�Q`V�҃���^��]����������hh�   h�f �|  ����t���   ��t��3��������U��hh�   h�f �I  ����t���   ��t]��]����U��M��U+u&�A+Bu�A+Bu�A+Bu�A+Bu�A+B]����������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���h�   h�   h�f �E��  �E��E��E�    �E�    �E�    ��  ����t���   ��t	�M�Q�Ѓ��UR�E�P��������]��U��E��u��MP�EPQ�s�����]��������������̋�3ɉ�H�H�H�U��V��~ W�}u0j j h8j��C������t
W���D���3��F��u_^]� �~ t3�9_��^]� ���H<�W�҃�3Ʌ����_�F   ^��]� �����V���F   ���H<�Q��3Ʌ����^���������������V��~ t�   ^Ã~ u3�^á��H<��AR�ЋN��Q���    �F    ����^����������U����u���H�]� ���J<�URP�A�Ѓ�]� ���������������U����u���H�]Ë��J<�URP�A�Ѓ�]�U����$V��u���H�1����J<�URP�A�Ѓ������Q�J`�E�SP�ы��B�Pp�M�QV�ҡ��H�A`�U�R�Ћ��Q�Jdj j��E�h{P�ы��Bj �M�Q�U�R�P$�M�Q�҅����H�Al�U�R���Ѓ�4��[t.���Q�u�B`V�Ћ��Q�Jl�E�P�у���^��]Ë��B�M��@,jQ�U�R�Ћ��Q�E�M�PQ�J0�E�P�ы��B�u�H`V�ы��B�Pp�M�VQ�ҡ��H�Al�U�R�Ѓ�(��^��]�U����$SV��u���H�1����J<�URP�A�Ѓ������Q�J`�E�P�ы��B�Pp�M�QV�ҡ��H�A`�U�R�Ћ��Q�Jdj j��E�h{P�ы��Bj �M�Q�U�R�P$�M�Q�҅����H�Al�U�R���Ѓ�4��t/���Q�u�B`V�Ћ��Q�Jl�E�P�у���^[��]Ë��B�M��@,jQ�U�R�Ћ��Q�E�M�PQ�J0�E�P�ы��B�P`�M�Q�ҡ��H�Adj j��U�h{R�Ћ��Qj �E�P�M�Q�J$�E�P�ы����B�Pl�M�Q���҃�@��t-���H�u�Q`V�ҡ��H�Al�U�R�Ѓ���^[��]Ë��Q�E��R,jP�M�Q�ҡ��H�U�E�RP�A0�U�R�Ћ��Q�u�B`V�Ћ��Q�Jp�E�VP�ы��B�Pl�M�Q�҃�(��^[��]�����������U����$SV��u���H�1����J<�URP�A�Ѓ������Q�J`�E�P�ы��B�Pp�M�QV�ҡ��H�A`�U�R�Ћ��Q�Jdj j��E�h{P�ы��Bj �M�Q�U�R�P$�M�Q�҅����H�Al�U�R���Ѓ�4��t/���Q�u�B`V�Ћ��Q�Jl�E�P�у���^[��]Ë��B�M��@,jQ�U�R�Ћ��Q�E�M�PQ�J0�E�P�ы��B�P`�M�Q�ҡ��H�Adj j��U�h{R�Ћ��Qj �E�P�M�Q�J$�E�P�ы����B�Pl�M�Q���҃�@��t-���H�u�Q`V�ҡ��H�Al�U�R�Ѓ���^[��]Ë��Q�E��R,jP�M�Q�ҡ��H�U�E�RP�A0�U�R�Ћ��Q�J`�E�P�ы��B�Pdj j��M�h{Q�ҡ��Hj �U�R�E�P�A$�U�R�Ћ��Q�Jl���E�P���у�@��t/���B�u�H`V�ы��B�Pl�M�Q�҃���^[��]á��H�U��I,jR�E�P�ы��B�M�U�QR�P0�M�Q�ҋu���E�P���������Q�Jl�E�P�у���^[��]���������U����$SV��u���H�1����J<�URP�A�Ѓ������Q�J`�E�P�ы��B�Pp�M�QV�ҡ��H�A`�U�R�Ћ��Q�Jdj j��E�h{P�ы��Bj �M�Q�U�R�P$�M�Q�҅����H�Al�U�R���Ѓ�4��t/���Q�u�B`V�Ћ��Q�Jl�E�P�у���^[��]Ë��B�M��@,jQ�U�R�Ћ��Q�E�M�PQ�J0�E�P�ы��B�P`�M�Q�ҡ��H�Adj j��U�h{R�Ћ��Qj �E�P�M�Q�J$�E�P�ы����B�Pl�M�Q���҃�@��t-���H�u�Q`V�ҡ��H�Al�U�R�Ѓ���^[��]Ë��Q�E��R,jP�M�Q�ҡ��H�U�E�RP�A0�U�R�Ћ��Q�J`�E�P�ы��B�Pdj j��M�h{Q�ҡ��Hj �U�R�E�P�A$�U�R�Ћ��Q�Jl���E�P���у�@��t/���B�u�H`V�ы��B�Pl�M�Q�҃���^[��]á��H�U��I,jR�E�P�ы��B�M�U�QR�P0�M�Q�҃�j h{�M��������Hj �U�R�E�P�A$�U�R�Ћ��Q�Jl���E�P���у����Q������H�U��I,jR�E�P�ы��B�M�U�QR�P0�M�Q�ҋu���E�P��襠�����Q�Jl�E�P�у���^[��]���������U����H<�A]����������������̡��H<�Q�����V��~ u>���t���Q<P�B�Ѓ��    W�~��t���j9��W�8�����F    _^��������U���V�E�P���Y����P���#����M���)9����^��]��̃= uK���t���Q<P�B�Ѓ��    ���tV����8��V�
8�����    ^������������U���8���H�A`S�U�V3�R�]��Ћ��Q�JdSj��E�h{P�ы��B<�P�M�Q�ҋ���H�Al�U�R�Ѓ�;�u^3�[��]�V�M�]���  �M�Q�U�R�M��(  ����   W�}�}���   �����   �U��ATR�Ћ�����tF���Q�J`�E�P���у��U�Rj�E�P���|������Qj WP�B �Ѓ��E���t�E� ��t���Q�Jl�E�P����у���t���B�Pl�M�Q����҃��}� u"�E�P�M�Q�M��[  ���7����E�_^[��]ËU��U�_�E�^[��]����������U��E����u��]�VP�M��  �EP�M�Q�M��E�    �E    ��  ����   �u�E���tB��t=��u[�����   �M�PHQ�ҋ��Qj VP�B �Ѓ���u-�   ^��]Ë����   �E�JTP��VP�V�������uӍUR�E�P�M��o  ���{���3�^��]�V��~ u>���t���Q<P�B�Ѓ��    W�~��t���:6��W�d5�����F    _^�������̋�� {���������{���������̅�t��j�����̡��P��l  ����P��x  ��U����P��p  ��V�E�P�ҋuP���z5���M��5����^��]� ��������̡��P��t  ��U����H��d  ]��������������U����H��  ]�������������̡��H��h  ��U����H��<  ]��������������U����H���  ]��������������U����H���  ]��������������U���EV���{t	V��Y������^]� �������������̸   � �������̸   @� �������̸   � �������̸   � ��������U����H�Q`V�uV�҃���^]� �3�� �����������3�� �����������U����   h�   ��@���j P��I  �M�Eh�   ��@���R�M��MPQjǅ`���    ����� ��]���U����   V�u��u3�^��]�h�   ��@���j P�uI  �M�U�Eh�   �M���@���Q�U��U��@����ERPj��`���ǅD������E�@��E����E�P��E����E�p��E�0��E�`������ ^��]�������������U���   SV�u(3ۉ]���u���H�Al�UR�Ѓ�^3�[��]Ë��Q�JW�EP3��у����'  �X,  �E���tq�UR�M��U2��Wh {�M�����P�M��>2���u�Wj��E�P�M�Q��\���R�_?�QR����P��x���P�4����P�M�Q�4����P���-  �E���t�E� �� t�M�����<2����t��x�������)2����t��\�������2����t�M̃���2����t���B�Pl�M�Q����҃���t�M���1���}� t"�E(�M$�U�P�EQ�MR�UPQR����������E�P�K+  ����M$�U�EVQ�Mj RPQ�����������B�Pl�MQ�҃���_^[��]�����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`�����������U������   �BXQ�Ѓ���u]� �����   �M�RQ�MQP�҃�]� U������   �BXQ�Ѓ���u]� �����   �M�R8Q�MQP�҃�]� U��EV��j ����Qj j P���   �ЉF����^]� ��Vj ��H����   j j R�Ѓ��F^�������������U��V��F��u^]� ���Q�MP�EP�Q���   P�у��F�   ^]� �U�����W��������Au���]��W���G��Au���]��E���z������A�  �E����������  ���0{������AuI������AuBV�[O  ���TO  �ȋ��ƙ����ʅ�u�u��E�^�]���E����������__��]�������������Au������=({��������Au>�����]������]������O�_�E��E�����������Au�����U��_�E�������������I �E��E����f  �]��E��]��E��U��${����t���E����������__��]���������__��]���������__��]����������������U��E��u�E�M�(�$�   ]� �����������U��EHV����   �$����   ^]á,@�,��uQ�EP�7�����=�*  }�����^]Ëu��t�j j h8j�,������t ����,��� ��tV���/���   ^]��     �   ^]ËM�UQR�����������H^]�^]�C����-,u.�e���� ���� ��t���/-��V�Y,�����     �   ^]Ã��^]Ë���6�=���|������U��E�M�UP��P�EjP�C}����]��������������̸   �����������U��V�u��t���u6�EjP�D}������u3�^]Ë��q~����t���t��U3�;P��I#�^]�������U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U��V�u�F��F�����������������]�E�_  �]�����E��������D�Ez��^�P�P�]��������]��E����������N�X�N^�X]�����������U�������P�P��P�P�P�P �P�P�P,�P(�P$�U�M��U��U��U����M��U�P�ɋU��U��U��P�U�H�U��U��M����U��H�M��ɉP�U�U��]��H�M��P�U��]��P$�U��H �M��H(�P,��]�������������U���`�M�A,V�I�A(�I ���I�A(�I�A�I,���I���A�I �A�I���I$���]���E��������Dz�u�؋��������^��]���W���]�A�I,�A�I(�A�I�A�I �A(�I �U��A,�I�]������I$�����I�����e��	���E�������]��A�I�U��A�I�]��A�I,�]��A(�I�U����e��I$�E�������������A�������������]��A�I�A�I �����	�����A�������E��e��I���E�ʍu��ɋ��]��E��e����]��E��e����]����������]��A$�I �A�I,�����]��A,�I�A$�I�����]��A�I�A �I�����]��A(�I�A$�I�����]��A$�I�A(�I�����]��A�I�A�I�   �����]��_^��]�����������U�������P�P��P�P�X�8{�@    �U��U��U��]�M��4{��M��U��U��P�]�U�P�U��H�M��H�P��]����������U��y t�U��������Au���B�A������Au�B�Y�B�A������Au�B�Y��A������z��Y�B�A������z�B�Y�B�A������z6�B�Y]� �E��Q�P�Q�@�A�Q�A��Q�A�Q�A   ]� ��������U����y ��   ��E�A�]��A�A�]��A�A�]��E���r�����]�U��E�����]�U�P�M��]��U��P�A� �]��A�`�]�U��A�M��`�E��P�]��M��H��]� ��E�U�V�u��U�U��]�M��P�p�E��P�p^��]� �������������̋�3ɉ�H�H�H�V����t	P�QG�����F�    ��t	P�;G�����F    �F    �F    ^��U��V��W��t	P�G�����F�    ��t	P��F�����}�F    �F    �F    ����   �? ��   �G����   3ɺ   ����j j h8���Q�qE�������t=� t?�G��t83ɺ   ����j j h8���Q�<E�����F��u�������_3�^]� �G��F�G��    Q�F�RP脉���F����t�N�W��QPR�h�����_�   ^]� ����������U��SV��3�W;�t	P��E�����F�;�t	P��E�����^�^�^9]��   �};���   3ɋǺ   ����SSh8���Q�iD�����;�t>9]tG�]��t@3ɋú   ����j j h8���Q�3D�����F��u�������_^3�[]� �^�13ɸ   �F�   ����j j h8���Q��C�����F��t���U��    PQR�~�L����E����t!�N�V��QRP�0�����_^�   []� �F�8_^�   []� 3���A�A�A���U��Q�A�`�
�@�b�	���B�a����]��E���]�������U���|��UV�U��q�<��M��E�    �,  S�]W���  ��Uԋ�UЋM�U̍@�<����}��x�@�E��B�@�����E��}����>��U����]��@�E��������]��@�E��E��E؋E�����E����]ȋEȉE�   ;��  �w����`  �w�����F�B��   �U�P��R�������]��B���]��B�U����]��E����E������E��M������]��E��E������E����������]��E��M؉U؋U����ɉU܋U�U���P��R���]��E��E��]��E��E��]��E��E��]�����]��B���]��B���]��E����E������E��M������]��E��E������E��ˋU��������]��E��M؉U؋U����ɉU܋U�U����R���]��E��E��]��E��E��]��E��E��]�����]��B���]��B�U����]��E����E������E��M������]��E��E������E����������]��E��M؉U؋U����ɉU܋U�U��P��R���]��E��E��]��E��E��]��E��E��]���������]��B���]��B�U����]��E����E������E��M������]��E��E������E����������]��E��M؉U؋U����ɉU܋U�U����]��E��E��]��E��E��]��E��E��]��������U�E��;���   �ۍ�+���@����������]��@���]��@�E����]��E����E������E��M������]��E��E������E����������]��E��M؉E؋E����ɉE܋E�E����]��E��E��]��E��E��]��E��E��]��g�������������������UȋE��UċU��]��M���S�M�Q�U�R�C��������ẺK$�ыP�S(�@�C,������z	�����]��U�E�������z	�����]���U��E�E������E�����   ��������z���]��������z	�����]���U��E�E�������zb�������C(�����C,���]��M��C$���C,�����]ċU��c$�K�S�]ȋEȉC�C�K(�C�K,���]��C�K,�C�K$�   �����������z���]��������z���]��E�E���������   �C,�����C(���]��M��C$�����]ċU��C$���C(�K�ʉS���]ȋEȉC�C(�K�C,�K���]��C,�K�C$�K�M����]ċU��C$�K�C(�K�K�S���]ȋEȉC �{�C(�����C,�������]��M��K$�C,���]ċU��c(�K�S�]ȋEȉC �C�K,�C �K(���]��M��C$�K �C,�K���]ċU��C(�K�C$�K�K�S���]ȋEȉC�M�SQ������U�   �����M������3�3�3���|'�y�����B�U�҉U�U�w����u�U�};�}�Q���U��U�9��E�Ƌu�E����@�����K��@�K���@�K$���]��C��C�@�K���C(�H���]��C��C�@�K ���C,�H�E��E��E����E��]ȋEȉE��E��D��@�����K��@�K���@�K$���]�� �K�C�@�K���C(�H���]�� �K�C�@�K ���C,�H�ẺE����]ԋEЋI���EċE�3��Eȅ���   �F���FU�;���@�E�����K�U���@�K���@�K$���]��C��C�@�K���C(�H���]��C��C�@�K ���@�E��K,���]��E����E������E��U��U��ʉU��E��U����E���E��E��E��E��ʉU��ʉE��������E������]�E�E��]��5����E�_[^��]� �������h0Ph_� ��������������������h0jh_� ���������uË@����U��V�u�> t/h0jh_� ��������t��U�M�@R�Ѓ��    ^]���U��Vh0jh_� ���i�������t�@��t�MQ����^]� 3�^]� �������U��Vh0jh_� ���)�������t�@��t�MQ����^]� 3�^]� �������U��Vh0jh_� �����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh0jh_� ����������t�@��t�MQ����^]� 3�^]� �������U��Vh0j h_� ���Y�������t�@ ��t�MQ����^]� 3�^]� �������U��Vh0j$h_� ����������t�@$��t�MQ����^]� 2�^]� �������Vh0j(h_� �����������t�@(��t��^��3�^������Vh0j,h_� ����������t�@,��t��^��3�^������U��Vh0j0h_� ���y�������t�@0��t�MQ����^]� 3�^]� �������U��Vh0j4h_� ���9�������t�@4��t�M�UQR����^]� ���^]� ��Vh0j8h_� �����������t�@8��t��^��3�^������U��Vh0j<h_� �����������t�@<��t�MQ����^]� ��������������U��Vh0j@h_� ����������t�@@��t�MQ����^]� ��������������U��Vh0jDh_� ���I�������t�@D��t�MQ����^]� 3�^]� �������U��Vh0jHh_� ���	�������t�@H��t�MQ����^]� ��������������Vh0jLh_� �����������t�@L��t��^��3�^������Vh0jPh_� ����������t�@P��t��^��^��������Vh0jTh_� ���l�������t�@T��t��^��^��������Vh0jXh_� ���<�������t�@X��t��^��^��������U��Vh0j\h_� ���	�������t�@\��t�M�UQR����^]� 3�^]� ���U��Vh0j`h_� �����������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh0jdh_� ����������t�@d��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh0jhh_� ���9�������t�@h��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh0jlh_� �����������t�@l��t�M�UQR����^]� 3�^]� ���U��Vh0jph_� ����������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh0jth_� ���i�������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh0jxh_� ���)�������t�@x��t�MQ����^]� 3�^]� �������U��Vh0j|h_� �����������t�@|��t�M�UQR����^]� 3�^]� ���U��Vh0h�   h_� ����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh0h�   h_� ���F�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U���X��A�U�V�U��]����z  S��E��EW����������O  ���������U�r�z�
�R;��4v���I�$��4����R����   �]��F�a�]��F�a�]���!�]��B�a�]��B�a�]��E����E������E����E����������]��E������E������������]��������]��E��E��]��E��E��]��E��   �]��F�a�]��F�a����]���!�]��B�a�]��B�a�]��E����E������E����E����������]��E������E������������]��������]��E��E��]��E��E��]��E��E��]����m������_[�u�E�PV���������^��]� U���$V��M�������F����   �6S�]W�u��E���$    ���������t[��%�����E�M܋���@��P�����F�@��R�M�������~���Q�M�������v;�t�v��P�M�������u����m��u�u�_[�M�UQR�M��v���^��]� ��������������̋Q3���|�	��t��~�    t@����u��3���������U��QV�u;��}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��|+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~#V�1�d$ ���   @u	�����t@����u�^���̋QV3���~�	�d$ ����ШtF����u��^���������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%���;��E���}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$����E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��2�H�[�o�������U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V����t	P�.�����F�    ��t	P�.�����F    �F    �F    ^��U��3�V���F�F�F�EP�D�����^]� �������������U��EVP���!�����^]� ����������U��SV��W3�;�t	P�.�����F�>;�t	P�.�����]�~�~�~;�to3ɋú   ����WWh8���Q�,�������tG�}��tI3ɋǺ   ����j j h8���Q�u,�����F��u���t	P�-�����    _^3�[]� �~_�^^�   []� �����������U��Q�A�E� ��~LS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U�����u�_^[�E��Ћ�]� ���������U��3�V��W�}��F�F�F�Gj;Gu2j������tY�����O�H�G��B�N_���   ^]� j�f�����t'�����W�Q��O�H��G�B�N�   _��^]� ��̡��H��   ��U����H��  V�u�R�Ѓ��    ^]����������̡��P��  Q�Ѓ�������������U����P�EPQ��  �у�]� ̡��H�������U����H�AV�u�R�Ѓ��    ^]��������������U����H�AV�u�R�Ѓ��    ^]��������������U����P��Vh�  Q���   �E�P�ы����   �Q8P�ҋ�����   ��U�R�Ѓ���^��]��������������̡��P�BQ�Ѓ����������������U����P�EPQ���   �у�]� �U����P�EP�EP�EP�EP�EPQ���   �у�]� �U����P�EP�EP�EP�EPQ�Jx�у�]� �������̡��P�B$Q��Y�U����P�EP�EP�EPQ�J�у�]� ������������U����P�EP�EP�EPQ�J �у�]� ������������U����P�EP�EP�EP�EPQ�J(�у�]� ��������U����P�EP�EPQ�J,�у�]� U����P�EP�EP�EPQ�J0�у�]� ������������U����P�EP�EP�EP�EPQ�J<�у�]� ��������U����P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U����P�EP�EP�EP�EPQ�J@�у�]� ��������U���V��H�QWV�ҋ����H�QV�ҋ��Q�M�RHQ�MQ�MQOWHPj j V�҃�(_^]� ���������������U����P�E P�EP�EP�EP�EP�EP�EPQ�JH�у� ]� ������������U����P�EP�EPQ�JX�у�]� U����P�EPQ�J\�у�]� ���̡��P�BlQ�Ѓ���������������̡��P�BpQ�Ѓ����������������U����P�EPQ�Jt�у�]� ����U����P�EP�EPQ���   �у�]� �������������U����P�E���   ��VP�EPQ�M�Q�ҋu�    �F    �����   j P�BV�Ћ����   �
�E�P�у� ��^��]� ������̡��P���   Q�Ѓ������������̡��H�������U����H�AV�u�R�Ѓ��    ^]��������������U����P�EP�EP�EP�EP�EP�EPQ�J�у�]� U����P�EPQ�J�у�]� ���̡��P�BQ��Y�U����P�EP�EPQ�J�у�]� U��VW�������M�U�x@�EPQR�������H ���_^]� �U��VW�������M�U�xD�EPQR���n����H ���_^]� �V���X����xH u3�^�W���F����΍xH�<����H �_^�����U��V���%����xL u3�^]� W�������M�U�xL�EPQR��������H ���_^]� �������������U���S�]VW���t.�M�視���������xL�E�P�������H ��ҍM������}��tZ���H�A`�U�R�Ћ��Q�Jp�E�WP�ы��B�Pl�M�Q�҃����Y����@@��t���QWP�Bp�Ѓ�_^[��]� ������U��VW���$����xH�EP�������H ���_^]� ���������U��VW��������M�U�xD�EP�EQRP��������H ���_^]� �������������U��V�������xP u
�����^]� W�������M�U�xP�EP�EQ�MR�UPQR���{����H ���_^]� ��������������U��V���U����xT u
�����^]� W���=����M�xT�EPQ���+����H ���_^]� ��������������U��V�������xX tW��������xX�EP��������H ���_^]� ������������U����MV3��E�PQ�u�u��u��u�u��  ����t.�E�;�t'���J�U�R�U�R�U�R�U�RP�Ax�Ѓ�^��]�3�^��]����������������h4Ph�f �������������������U��h4jh�f �l�������t
�@��t]�����]�������U��Vh4jh�f �;���������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�����E�NP�у�4�M��������^]ÍM�������^]��U��h4jh�f ���������t
�@��t]��3�]��������U��h4jh�f ��������t�x t�P]��3�]Ë�U���V�u��u�W?  �@�E��&?  ���E�F�}� �E�u�E�H�����   �� ��   S�]W�   ;�s��uS�9  Y��u�   �F�Xt}��u�]��}��t8  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPW�u�j ��7  ��$��u������E�t	�M����_[^�Ë�U��V�T>  �@�u��!>  jh   �F�>  YY�F��th   �7  P�v�  ���F   ��7  �f �F��^]Ë�Whl����p��uV�@V��  �����Y|�^��_�hl��p��}V�@V�  �����Y|�^Ë�U��E��V��}k�@P�  Y��^]� ���}k�@P�  YË�U���u��1  Y��t]�2?  ]ËI������t�j���Ë�U��V��������EtV���Y��^]� ��U��E���t�|�����t�j���]Ë�U��Qj �M��@���h�������%� Y�M��N����á�Ë�U��=� uh������  Y�E��]�j�Qj�?  j �M�������}�e� �w��GN���8 t��������t�j�����w��w�x  �M��Y�M�������?  Ë�U��Qj �M�������ȋ j�����������u�M������Ë�U��=� uh������Yj����Y��t����M�H�3���]Ë�U��E�xP v�xTr�@@���@Pj �YM  YY]�j�tj�>  ��u��F   3��E��F�F�F�EhP{�N�L{�F�hZ�����>  � j��j�D>  ��u��L{V�E�   ����Yj j�N�}A���Pu�}>  Ë�U��V�������EtV����Y��^]� j��j��=  ������u{P�M��2�����!u�����uXj4����Y�ȉM��E���t
V�������3�V�E� ������N�F?   �$T{�aQ���Ή5�����������M���M����������=  Ë�U��E�xVWr�p��pj j ��K  YY��u��r�}P�O<��P����tVj ��K  YY��u�P{P�OX��P��_^]Ë�U��VW���w ��vW�u�V�6����u�_^]� ��U��V�uWj ��������F��t�8P���Y�ǅ�u�F �f ��t�8P���Y�ǅ�u�f  _^]Ë�U��V�u�~ v�F���F�� V����Y�N$��tj�_&��^]Ë�Vj���`��P��2  YY��^Ë�V���6�0  �6���YY^��1�.  Y��1�5  YË�U���V�u��u��8  �@�E���8  ���E�F�}� �E�u�E�H�����   �� ��   S�]��   s!��uS�63  Y��u�   �F�X��   ��u�]��}��2  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPh   �u�j �g1  ��$��u������E�t	�M����[^�Ë�U��V�u���T���`{��^]� �`{�T����U��V���`{�lT���EtV���Y��^]� jD��j�:  hh{�M��V���e� �E�P�M��T��h���E�P�X  �jD��j�f:  hx{�M��gV���e� �E�P�M��P���h@��E�P�   ̋�U��V�u���]���`{��^]� ��U��USVW�ڋ�����   ��@t����t��3Ɂ�;���3�A;�t���{@��u��������{ u3��^��t%��t �uh�{�u��I  ����t	P��#  Y���u����V�u�I  ������t���tjj V�h"  ����tV�ŋ�_^[]Ë�U���  �p�3ŉE��Eh  Ph  ������Pj ��L  ����t3���u�������uP��������M�3��  �Ë�U���u� p]Ë�U���u�$p]Ë�U���u�(p]Ë�U���u�,p]Ë�U�����u]�7  �MH����0]����0@����t��,����
r������������̋L$WSV��|$��to�q��tU���L$���:�t��t���:�t
��u�^[_3�Ê��:�u�~��a��t(���:�u��A��t�f���:�t��3�^[_����K  �G�^[_Ë�^[_Ë�U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$����U��QQSVWd�5    �u��E�:�j �u�u��u��~ �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�W  �� �E�_^[�E���]Ë�U��V��u�N3��  j V�v�vj �u�v�u�kW  �� ^]Ë�U���8S�}#  u�w��M�3�@�   �e� �Eܣ��p��M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E��Z  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M�  �E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u�5V  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����-���u�	]  �M�N��k���M9H};H~���u	�M�]�u�} }ʋEF�0�E�;_w;�v��\  ��k�E�_^[�Ë�U��EV�u��Y  ���   �F�Y  ���   ��^]Ë�U����X  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V��X  �u;��   u�X  �N���   ^]��X  ���   �	�H;�t���x u�^]�\  �N�H�ҋ�U����p��e� �M�3��M�E��E�E�E@�E���M��E�d�    �E�E�d�    �uQ�u�\  �ȋE�d�    ����;p�u���A\  ��Q�$|�9]  YË�U��V��������EtV����Y��^]� ��U��E��	Q��	P�]  ��Y�Y@]� ��U��E��t���8��  uP�  Y]Ë�U��EV���F ��uc�W  �F�Hl��Hh�N�;x�t����Hpu�6  ��F;��t�F����Hpu�_  �F�F�@pu�Hp�F�
���@�F��^]� ��U����p�3ŉE�S3�V;�u�xd  j^SSSSS�0�  ���5  �uW��c  YY;Er��ЋU��H;�u ��8t�<a|<z, �A8u�3���   j�p�   SSj�WVQR�(  �ȃ�$�M�;�u��c  � *   ��c  � �   9Ms���c  j"�^���;�~Ej�3�X���r9�A=   w�d  ��;�t� ��  �P��   Y;�t	� ��  ���M�E���]�9]�u�~c  �    냋U�j�pQ�u�j�WV�pR�(  ��$��t�u��uW��   ������<c  j*Y����u������Y�ƍe�^[�M�3��}����Ë�U���W�u�M�������}�E�P�u�_����}� YY_t�M��ap��Ë�U��j �u�u������]Ë�U��S3�9�uA�E;�u�b  SSSSS�    �  ��3��/��8t)�
��a|
��z�� �
B8u��Sj��u�X����E��[]Ë�U��MS3�VW;�t�};�w�Kb  j^�0SSSSS�S  �����0�u;�u��ڋъ�BF:�tOu�;�u��b  j"Y�����3�_^[]������̋T$�L$��ti3��D$��u��   r�=�* t�b  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�ø9@� ��� 7���6��7��v6�����?���6� ��5�$��5Ë�U�������n  �} �`t�#n  ��]��̃=�* �fq  ���\$�D$%�  =�  u�<$f�$f��f���d$�5q  � �~D$f(P|f(�f(�fs�4f~�fT�|f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$��m  ���D$��~D$f��f(�f��=�  |!=2  �fT@|�\�f�L$�D$����f�p|fVp|fT`|f�\$�D$���������������̃=�* �q  ���\$�D$%�  =�  u�<$f�$f��f���d$��p  � �~D$f(�|f(�f(�fs�4f~�fT�|f��f�ʩ   tL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$��l  ���D$��~D$f��f(�f��=�  |%=2  �fT�|�X�f�L$�D$���|�f��|fT�|f�\$�D$����U��WV�u�M�}�����;�v;���  ��   r�=�* tWV����;�^_u^_]�q  ��   u������r*��$�$���Ǻ   ��r����$�8��$�4���$����H�t���#ъ��F�G�F���G������r���$�$��I #ъ��F���G������r���$�$��#ъ���������r���$�$��I �� ������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�$���4�<�H�\��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$�p��I �Ǻ   ��r��+��$����$�������� ��F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I t�|��������������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�������������U��WV�u�M�}�����;�v;���  ��   r�=�* tWV����;�^_u^_]�m  ��   u������r*��$�����Ǻ   ��r����$����$�����$�(�������#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I ��x�p�h�`�X�P�H��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�0������$����I �Ǻ   ��r��+��$�4��$�0��D�h����F#шG��������r�����$�0��I �F#шG�F���G������r�����$�0���F#шG�F�G�F���G�������V�������$�0��I �����������'��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�0���@�H�X�l��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̃=�* t-U�������$�,$�Ã=�* t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$�Ë��` �` � �|Ë�U��S�]VW����|���t&P�#  ��FV�,  YY�G��t�3VP�l�������g �G   ��_^[]� ��U��S�]V����|�C�F���CWt1��t'P�W#  ��GW��  YY�F��t�sWP�������	�f ��F_��^[]� �y ��|t	�q��  YËA��u��|Ë�U��V�EP��������|��^]� ��U��V�u���R�����|��^]� ��|������U��V�������EtV�B��Y��^]� ��U��V����|�c����EtV���Y��^]� ��U��V�uW3�;�u3��e9}u�U  j^�0WWWWW�  �����E9}t9urV�u�u���������uW�u�X�����9}t�9us�@U  j"Y����jX_^]������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[Ë�U��EVW3�;�tG9}u�cT  j^�0WWWWW�k  �����)9}t�9Es�>T  j"Y�����P�u�u�������3�_^]Ë�U��E�d]Ë�U���(  �p�3ŉE������� SjL������j P�������������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������Dpj ���@p��(���P�<p��u��uj�f  Yh ��8pP�4p�M�3�[�M����Ë�U���5d�C  Y��t]��j�Wf  Y]����3�PPPPP�������Ë�U��� �EVWjY�}�}��E��E_�E�^��t� t�E� @��E�P�u��u��u��Hp�� jh���	s  �u��tu�=|*uCj��g  Y�e� V�!h  Y�E��t	VP�Bh  YY�E������   �}� u7�u�
j��f  Y�Vj �5�Pp��u��Q  ���LpP�Q  �Y��r  �jh���{r  3��}�3��u;���;�u �Q  �    WWWWW����������   V�u  Y�}��F@uwV�y  Y���t���t�����ȃ����@����A$u)���t���t���������@����@$�t�*Q  �    WWWWW�1������M��9}�u�Nx
��A��V�Pu  Y�E��E������   �E���q  ËuV��t  Y�jh���wq  3��}�3��u;���;�u �P  �    WWWWW����������   V�	t  Y�}��F@uwV�x  Y���t���t�����ȃ����@����A$u)���t���t���������@����@$�t�&P  �    WWWWW�-������M��9}�u!�Nx��E�����V�u�Dx  YY�E��E������   �E���p  ËuV�s  YË�U��V�u�F@WuyV��w  Y�����t���t�ȃ��������@����A$u&���t���t�ȃ������@����@$�t�ZO  3�WWWWW�    �_���������JS�]���t=�F�u��y2�u.3�9~uV��x  Y�;Fu9~u@���F@�t8t@����[_^]È�F�F�����F��%�   ��jh��zo  3�3�9u��;�u�N  �    VVVVV�����������+�u�r  Y�u��u�u�����YY�E��E������	   �E��do  ��u�Tr  YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�Vv  YP�a  ��;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV��u  P��  Y��Y��3�^]�jh(��Xn  3��}�}�j�Pc  Y�}�3��u�;5`*��   �@��98t^� �@�tVPV�%q  YY3�B�U��@���H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u�@�4�V�.q  YY��E������   �}�E�t�E���m  �j�a  Y�jhP��~m  3�9uu	V����Y�'�u�1p  Y�u��u����Y�E��E������	   �E��m  ��u�wp  Y�j�����Y�jhp��"m  3ۉ]�3��u;���;�u �\L  �    SSSSS�c���������   �E��t	;�t��@u�;�t��@u�}�G�=���v뷋}����uV�o  Y�]�V����V��~  YY�f�����N�Et���Fj_�-�E;�u W�b  Y;�u�d�M����N  �	��   �N�~�F��^�E������	   �E��l  ��u�po  YË�U���SVW3�9}t$9}t�u;�u�_K  WWWWW�    �f�����3�_^[�ËM;�tڃ��3��u9Ew͋}�}�F  �M��}��t�F�E���E�   ����   �N��  t/�F��t(��   ��;�r��W�u��6�-���)~>��+�}��O;]�rO��tV�S���Y��u}�}� ��t	3ҋ��u�+�W�u�V�r  YP��{  �����ta��;�w��M�+�;�rP�}��)�E�� VP�r  YY���t)�E��FK�E����E�   ���A����E������N ��+�3��u������N �E���jh����j  3�9ut)9ut$3�9u��;�u ��I  �    VVVVV�������3���j  ��u�Mm  Y�u��u�u�u�u�=������E��E������   �E����u�m  YË�U��W3�9}u�I  WWWWW�    ����������AV�u;�u�gI  WWWWW�    �n����������u�  Y�ȉ#ʃ���V;�t3�^_]Ë�U��V�u�F��u�I  �    ����g���}�FuV�	�  E�e YV�����FY��y����F��t�t�   u�F   �u�uV��p  YP��  3Ƀ������I��^]�jh���Hi  3�3�9u��;�u�H  �    VVVVV����������>�};�t
��t��u��u��k  Y�u�W�u�u�������E��E������	   �E��i  ��u�l  YË�U��V3�9uu�H  VVVVV�    �����������E;�t�V�p�0�u�&�  ��^]Ë�U��SV�uW3����;�u��G  WWWWW�    ���������B�F�t7V�:���V���z  V�o  P軂  ����}�����F;�t
P����Y�~�~��_^[]�jh���h  �M��3��u3�;���;�u�@G  �    WWWWW�G����������F@t�~�E��
h  �V�j  Y�}�V�*���Y�E��E������   �ՋuV��j  YË�U��Q�e� S�]��u3��   W��ru�{���vn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9}�r��?�@��I��F�@��I��<�@��I��2�@��I��(�M�E����t:u@A�E�9]�r�3�_[��� �	+����U���u�Tp��u�Lp�3���tP�)F  Y���]�3�]Ë�U��� WV�  3�Y;�u��E  WWWWW�    �����������49}t޹����E�I   �u�u��M�;�w�E��u�E��u�uP�U��_�Ë�U��V�u�EPj �uh p�z�����^]Ë�U��j
j �u��  ��]Ë�U��EVW��u|P��X  Y��u3��  �l9  ��u��X  ���{�  �\p��*�4�  �l�j  ��}��5  ���_�  ��| �ޖ  ��|j 诔  Y��u�h�   �l  ��3�;�u19=h~��h9=�u�>�  9}u{�wl  �5  �\X  �j��uY�>5  h  j�W  ��YY;��6���V�5T��5��4  Y�Ѕ�tWV�w5  YY�Xp�N���V�����Y�������uW��7  Y3�@_^]� jh����d  ����]3�@�E��u9h��   �e� ;�t��u.�$}��tWVS�ЉE�}� ��   WVS�r����E����   WVS謝���E��u$��u WPS蘝��Wj S�B����$}��tWj S�Ѕ�t��u&WVS�"�����u!E�}� t�$}��tWVS�ЉE��E������E���E��	PQ�G�  YYËe��E�����3�� d  Ë�U��}u�B�  �u�M�U�����Y]� jh��c  �e� �u;5l*w"j�X  Y�e� V�`  Y�E��E������	   �E��c  �j�W  YË�U��V�u�����   SW�=`p�= u���  j�G�  h�   ��  YY�|*��u��t���3�@P���uV�S���Y��u��uF�����Vj �5�׋؅�u.j^9�t�u�ל  Y��t�u�{����B  �0�B  �0_��[�V谜  Y��A  �    3�^]Ë�U��� S3�9]u��A  SSSSS�    �����������N�E;�t�V�u�E��u�E��u�E�P�E�����E�B   ��  ���M��x�E����E�PS��i  YY��^[�Ë�U���uj �u�u�m�����]��������������̀�@s�� s����Ë������������Ë�U��QSVW�5(�M1  �5$���}��=1  ��YY;���   ��+ߍC��rwW芩  ���CY;�sH�   ;�s���;�rP�u���  YY��u�G;�r@P�u���  YY��t1��P�4��X0  Y�(�u�J0  ���V�?0  Y�$�EY�3�_^[�Ë�Vjj �;  ��V�0  ���(�$��ujX^Ã& 3�^�jh0���`  規  �e� �u�����Y�E��E������	   �E���`  �腏  Ë�U���u���������YH]�̺��顩  �����  �Ƀ=`t����d�  �����z�����������������̃��$譻  �   ��ÍT$�X�  R��<$�D$tQf�<$t��  �   �u���=\ ���  �   ��逻  �  �u,��� u%�|$ u����  �"��� u�|$ u�%   �t����-��   �=\ �&�  �   ���/�  ZË�U����p�3ŉE�SV3�W��9|u8SS3�GWh(}h   S�pp��t�=|��Lp��xu
�|   9]~"�M�EI8t@;�u�����E+�H;E}@�E�|����  ;���  ����  �]�9] u��@�E �5lp3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�L>  ��;�t� ��  �P�(���Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5ppSSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�=  ��;�tj���  ���P�f���Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�pp��t"SS9]uSS��u�u�u�VS�u �hp�E�V����Y�u������E�Y�Y  �]�]�9]u��@�E9] u��@�E �u蠹  Y�E���u3��!  ;E ��   SS�MQ�uP�u 边  ���E�;�tԋ5dpSS�uP�u�u�։E�;�u3��   ~=���w8��=   w�w<  ��;�t����  ���P�P���Y;�t	� ��  �����3�;�t��u�SW��������u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u���  ���u������#u�W�_���Y��u�u�u�u�u�u�dp��9]�t	�u�����Y�E�;�t9EtP�����Y�ƍe�_^[�M�3������Ë�U����u�M������u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap����-  �ȋAl;x�t����Qpu�  ���   Ë�U����u�M������E����   ~�E�Pj�u迹  ������   �M�H���}� t�M��ap��Ë�U��=� u�E�h��A��]�j �u����YY]Ë�U����u�M��-����E����   ~�E�Pj�u�@�  ������   �M�H���}� t�M��ap��Ë�U��=� u�E�h��A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u���  ������   �M�H���}� t�M��ap��Ë�U��=� u�E�h��A��]�j �u����YY]Ë�U����u�M��/����E����   ~�E�Ph�   �u�?�  ������   �M�H%�   �}� t�M��ap��Ë�U��=� u�E�h��A%�   ]�j �u�~���YY]Ë�U����u�M������E����   ~�E�Pj�u輷  ������   �M�H���}� t�M��ap��Ë�U��=� u�E�h��A��]�j �u����YY]Ë�U���L�p�3ŉE�S3�V�uW�]ԉ]�]��]؉]܉u��]�9^�  �F9u P�F0h  P�E�SP��  ������  j�  j��  W�E��  jW�E��  jW�E��  jh  �E��  ��$�E�9]��|  9]��s  ;��k  9]��b  9]��Y  �Eԉ3��M܈@=   |�E�P�v�tp���/  �}��%  �E���E�~-8]�t(�E�:�t�x�����M�� �G;�~�@@8X�uۋE�SS�v   Ph   �u܉E�jS聸  �� ����  �M��E�S�v��   W���   QW@Ph   �vS������$����  �E�S�v�   WP�E�W@Ph   �vS�U�����$���`  �E�}����   3҃}�f��U؉Mč��   �_�Z��M����   �MȈ~S8]�tN�M�M�:�tB�I���;ʉM�'��H   ��M��E� �  f�AA�M̋M��	9M�~�M�AA�M�8Y�u�h�   ��   QP�M���j��   PW�>����E�j��   QP�,������   ��$;�tKP�p��u@���   -�   P�F������   ��   +�P�3������   +�P�%������   �������E��    ���   �E����   �Eĉ��   �E����   �Eȉ��   �EЉ��   �u������Y���m�u�������u������u������u�����3ۃ�C�ˍ��   �;�tP�p����   ǆ�   0~ǆ�   ��ǆ�   8�ǆ�      3��M�_^3�[�������8'  �ȋAl;x�t����Qpu�Q  �@��'  �ȋAl;x�t����Qpu�+  ��Ë�U��VW3��u������Y��u'9�vV�p���  ;�v��������uʋ�_^]Ë�U��VW3�j �u�u�յ  ������u'9�vV�p���  ;�v��������uË�_^]Ë�U��VW3��u�u詶  ��YY��u,9Et'9�vV�p���  ;�v��������u���_^]Ë�U��VW3��u�u�u�s�  ������u,9Et'9�vV�p���  ;�v��������u���_^]��̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U���(  �p�3ŉE�� �Vtj
�E�  Y�O�  ��tj�Q�  Y� ���   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P���������������(�����0���j ǅ����  @��������,����@p��(���P�<pj��  �Pd�5    �D$+d$SVW�(��p�3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(��p�3�P�e��u��E������E�d�    ËM�d�    Y__^[��]QË�U��SV�u���   3�W;�to=@th���   ;�t^9uZ���   ;�t9uP�t������   ��  YY���   ;�t9uP�S������   �a�  YY���   �;������   �0���YY���   ;�tD9u@���   -�   P�������   ��   +�P��������   +�P��������   ����������   �=�t9��   uP�λ  �7����YY�~P�E   ����t�;�t9uP����Y9_�t�G;�t9uP����Y���Mu�V�q���Y_^[]Ë�U��SV�5pW�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{���t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5pW�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{���t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�V���t��t;�tWj6Y���  P����Y_^Å�t7��t3V�0;�t(W�8����Y��tV�����> Yu����tV�3���Y��^�3��jhP���N  �   ����Fpt"�~l t�   �pl��uj �}  Y����N  �j�C  Y�e� �Fl�=x��i����E��E������   ��j�B  Y�u�áx��H� �H����   �|����   �8���   �p���   �����   �tË�U��SW�}3�;�~,V�u���6�u�u�q�  ����tSSSSS�7�����Ou�^_[]Ë�U��SVW�}h�   3�SW�*����u�����u3���   <.u4�F8t-jP���   jP���  ����tSSSSS����������   ��h@�V�]�a�  ;��   �} �<0�u��@��   ��.��   PVj@�u�;�}u��@sw��_trP�EVj@��@��}u`��s[��t��,uRP�EVj��P�:�  ����t3�PPPPP�:�������,�'����������E�wh@�V輿  ��YY�X������_^[]Ë�U��SV�uV�u�u������3ۅ�tSSSSS��������F@8tPhD�j�u�u�Q��������   8^[tPh(yj�u�u�/�����]Ë�U���S3�ChU  �]��!���Y�E���U  W�x� ��]��^�CH�0�E�hL��5��jhQ  W������E���E��E���hH�hQ  W�K�  ����t3�PPPPP�������sX�E��0�F#  YY��t�e� �E��E��E����0�CH�0�E�E�hL��0jhQ  W�Z������}���|��}� uI�FP�p��tP�Ӆ�u	�vP�B���Y�FT��tP�Ӆ�u	�vT�+���Y�E�fT �fL �FP�~H���N�u������FP�=p3�Y;�tP�ׅ�u	�vP�����Y�FT;�tP�ׅ�u	�vT�����Y�Fh�^T�^L�^P�^H_[�Ë�U���   �p�3ŉE��ESV�uW�}��d����E��\�����`����s  �   �H(��T����H,�X �   ��X�����h�������  ��d��� ��  �} ��  �>CuW�~ uQhT{�u��d����%�����3���tVVVVV�i�����;�t3�f�f�Gf�G��`���;�t�0��d����G  V������   Y��P���;�s,V��h����c!  YY����   V��X����M!  YY����   ��L��� ��l���VP����YY����   ��l���PSP�-�  ������   �C��T������l���PW��h����������> t
��P���;�r��L�����r@PVW��X����g�  ����t3�VVVVV�g������3�9�\���tjS��\���������9�`���tj��T�����`�����������h����u��d�����������tVVVVV��������h����3��M�_^3�[�]����Ë�U����  �p�3ŉE�SW���_  �u����h���P��P���Ph�   ��x���PS���  ��������u3��  �E���0�sH��x���P��  YY���x  ��x���P�:�����P��t��������YY��p�����t��CH�M��\����D���k���l���� ��X����1jP��d�����<���P�s����F��x���Q��t�����L�����p��������QP��������t3�PPPPP���������p�����l������CH��P����j��P���P��d����������}��   ��h�����t��� �F�G$�O ��d����ǋV;t6���t������d�����D����P�H��D�������t�����d���|��"��t�����t�ǋ��P�W���d����H��t���uhj�v��x����vPjh��jj �~�  �� ��t93���  f!�Ex���@��r�h�   �5$���x���P��  �����@�G��g �F��G���   �}u	��h����F�Ek�V����Y��t1��\�����p����CH������X���Y��l������L����F������\�����t-�E�����<0�7�p��u�7������sT�����cL YY�M��p��������    �1�CH�M�_3�[�[����Ë�U���   �p�3ŉE��ESV3ۋ�W��h���;�t;�tP�����Y��  ���D0H��  ǅp���   ��t���;���  �9L�0  �yC�&  �y_�  ��hP�W�6�  ��YY����   +ǉ�p�����   �;;��   ǅl���   ������p���PW�6�D�������u�6�����Y9�p���t��l���������~�ChH�S菷  ��3�YY;�u	�;;��   ��l���QWS��x���h�   P覷  ����tVVVVV��������l�����h�����x���Ƅ=x��� ����Y��t��t�����? t
G�? � ���3�9�t�����   ��h����u3��vSSSh�   ��x���PQ�"�����;�tZ�~H��t3�7��x���P�f  YY��tS��x����%���Y��u!�p������t���C����~�3�9�p���u9�t���t�D����M�_^3�[�@�����jhp��~C  3ۉ]��}v��"  �    SSSSS�������3��,  �%  ���u��Q����Np�]�jh�   �\���YY���}�;���   j�#8  Y�E�   �Nl�������]��   �u�M���P���Y�E�;���   9]th���u�_  YY��t
��   j��7  Y�E�   �^l���|���W����Y�Fpu2���u)�;�x��Z���j�x���Ph�������������e� �   �-�}܋u�3�j�6  YËu�j�v6  Y��W�N���W�p���YY�E������   �E��hB  Ëu�fp��jh���B  3��u�3��];���;�u�H!  �    VVVVV�O�����3��{3��};���;�t�3�f97��;�t����  �E;�u�!  �    �ɉu�f93u ��   �    j��E�Php����  ���P�uWS���  ���E��E������	   �E��A  ��u�D  YË�U���SV�u3ۉ]�;�t9]u3��{  v3�f�W�};�u�p   SSSSS�    �w������<  �u�M��/����E�;���   9XuH9]v�M��9f�f�8tAFF�M�;Mr�8]�t�E�`p��E���   8]�t�E�`p�����   �uVj�W�=lpj	�p��;���   �Lp��zt��  � *   3�f��   �E�u�E�;�t'��M�:�t�M���QP���  YY��tF8t!F9]�u��u+u�u�E�V�uj�p��;�uT�e  �M� *   3�f��-9Xu	W����Y�1SSj�Wj	�p�lp;�u�.  � *   8]�t�E�`p�����H8]�t�M�ap�_^[�Ë�U���SV�u3ۉ]�;�u9]t*�9]w��  j^SSSSS�0�����������   3�f�W�};�t��u�M�荹���E;Ev�E=���v	�  j�P�M�QP�uV����������u;�t3�f��l  � 8]�tk�M�ap��b@;�tH;Ev<�}�t,3�f��B  j"^SSSSS�0�J�����8]�t�E�`p����&�E�E�P   3�f�LF�;�t�8]�t�E�`p��E�_^[�Ë�U��j �u�u�u�u�u�������]�����������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[Ë�U��V�EP��������\���^]� �\��u�����U��V���\��b����EtV����Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR�  YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =MOC�t=csm�u+�  ���    ��  �  ���    ~�  �   �3�]�jh���<  �}�]��   �s��s�u��\  �   � �e� ;ute���~;w|��  �����Oȋ1�u��E�   �y t�sh  S�O�t��  �e� ��u��-���YËe�e� �}�]�u��u���E������   ;ut�a  �s�8<  Ë]�u��  ���    ~�  �   �Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�q  3�A��  ���3��jh���;  �M��t*�9csm�u"�A��t�@��t�e� P�q�V����E������;  �3�8E��Ëe��R  ̋�U��M�V�uƃy |�Q�I�42���^]Ë�U�����u
�c  �  �e� �? �E� ~SSV�E�@�@��p��~3�E����E�M�q�P�GE�P�_�������u
K�������E��E��E�;|�^[�E���j�k�t����X  ���    t��  �e� �  �M���|  �3  �Mj j ���   ������j,hh��>:  �ً}�u�]�e� �G��E��v�E�P�̲��YY�E���  ���   �E���  ���   �E���  ���   ��  �M���   �e� 3�@�E�E��u�uS�uW�������E�e� �o�E������Ëe��  ��   �u�}�~�   �O��O�^�e� �E�;Fsk�ËP;�~@;H;�F�L�QVj W�������e� �e� �u�E������E    �   �E��u9  ��E�맋}�u�E܉G��u�����Y��
  �Mԉ��   ��
  �MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v蚱��Y��t�uV�%���YY�jh���8  3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w�2�  YY����   SV�!�  YY����   �G��M��QP�����YY���   �}�E�p�tH���  YY����   SV���  YY����   �w�E�pV����������   ���t|��W�9Wu8��  YY��taSV��  YY��tT�w��W�E�p�_���YYPV襻�����9�e�  YY��t)SV�X�  YY��t�w�J�  Y��t�j X��@�E���  �E������E��3�@Ëe��Q  3��u7  �jh���#7  �E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS�Ѭ����FP�w����YYP�vS跬���E�������6  �3�@Ëe��  ̋�U��} t�uSV�u�V������}  �uuV��u �u����7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP�����]Ë�U��QQV�u�>  ���   W��  ���    t?��  ���   �z  9t+�>MOC�t#�u$�u �u�u�u�uV虬��������   �}� u�"  �u�E�P�E�PV�u W�������E���;E�s[S;7|G;wB�G�O����H��t�y u*�X��@u"�u$�u�u j �u�u�u�u�����u���E��E���;E�r�[_^�Ë�U���,�MS�]�C=�   VW�E� �I��I����M�|;�|�h
  �u�csm�9>��  �~� ��  �F;�t=!�t="���   �~ ��   �  ���    ��  �  ���   �u�q  ���   jV�E�l�  YY��u��	  9>u&�~u �F;�t=!�t="�u�~ u�	  �&  ���    t|�  ���   �  �u3����   ����Y��uO3�9~�G�Lh4��������uF��;7|��	  j�u�d���YYhd��M��7���h���E�P�r����u�csm�9>��  �~�~  �F;�t=!�t="��e  �}� ��   �E�P�E�P�u��u W蹫�������E�;E���   �E�9��   ;G|�G�E�G�E��~l�F�@�X� �E��~#�v�P�u�E����������u�M��9E���M�E��}� ��(�u$�]��u �E��u��u�u�uV�u�K����u���E����]����}�} t
jV�:���YY�}� ��   �%���=!���   �����   V����Y����   �_  �Z  �U  ���   �J  �}$ �M���   Vu�u��u$�^����uj�V�u�u�������v�����]�{ v&�} �)����u$�u �u�S�u�u�uV������� ��  ���    t�_  _^[�Ë�U��V�u���{����\���^]� ��U��SVW�  ��   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������� 3�@_^[]Ë�U��V�5X��5�p�օ�t!�T����tP�5X����Ѕ�t���  �'���V�xp��uV��^  Y��tht�P�|p��t�u�ЉE�E^]�j ����YË�U��V�5X��5�p�օ�t!�T����tP�5X����Ѕ�t���  �'���V�xp��uV�V^  Y��th��P�|p��t�u�ЉE�E^]���p� ��V�5X���p����u�5��e���Y��V�5X���p��^áT����tP�5��;���Y�ЃT���X����tP��p�X���`#  jh��~/  ���V�xp��uV�]  Y�E�u�F\�3�G�~��t$ht�P�|p�Ӊ��  h���u��Ӊ��  �~pƆ�   CƆK  C�Fhp�j�$  Y�e� �vh�p�E������>   j��#  Y�}��E�Fl��u�x��Fl�vl�N���Y�E������   �/  �3�G�uj��"  Y�j��"  YË�VW�Lp�5T��������Ћ���uNh  j������YY��t:V�5T��5������Y�Ѕ�tj V�����YY�Xp�N���	V�$���Y3�W��p_��^Ë�V��������uj�t\  Y��^�jh0��.  �u����   �F$��tP�׺��Y�F,��tP�ɺ��Y�F4��tP軺��Y�F<��tP譺��Y�F@��tP蟺��Y�FD��tP葺��Y�FH��tP胺��Y�F\=�tP�r���Yj�"  Y�e� �~h��tW�p��u��p�tW�E���Y�E������W   j�M"  Y�E�   �~l��t#W�@���Y;=x�t����t�? uW�L���Y�E������   V����Y�A-  � �uj�!  YËuj�!  YË�U��=T��tK�} u'V�5X��5�p�օ�t�5T��5X����ЉE^j �5T��5�����Y���u�x����X����t	j P��p]Ë�VW���V�xp��uV�Z  Y�����^  �5|phІW��hĆW����h��W����h��W���փ=� �5�p��t�=� t�=� t��u$��p����p��$�5�����p�X������   �5�P�օ���   �\  �5������5��������5��������5����u���������  ��teh�%�5������Y�УT����tHh  j�V�����YY��t4V�5T��5�����Y�Ѕ�tj V�y���YY�Xp�N��3�@��$���3�_^�jhX���*  �����@x��t�e� ���3�@Ëe��E������V�����*  ��~����@|��t������jhx��*  �5�����Y��t�e� ���3�@Ëe��E������}����h")�g���Y������������U���SQ�E���E��EU�u�M�m��%�  VW��_^��]�MU���   u�   Q��  ]Y[�� ��U���(  ���������5��=�f��f��f��f��f�%�f�-�����E ���E���E����������  ������	 ���   �p��������t��������Dp��j�  Yj �@ph܆�<p�=� uj��  Yh	 ��8pP�4p��jh����(  j��  Y�e� �u�N��t/�����E��t9u,�H�JP螵��Y�v蕵��Y�f �E������
   ��(  Ë���j�  Y��������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP����3��ȋ��~�~�~����~����p����F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �p�3ŉE�SW������P�v�tp�   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R�?�����C�C��u�j �v�������vPW������Pjj 菇  3�S�v������WPW������PW�vS������DS�v������WPW������Ph   �vS�~�����$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[耟����jh���%  ����������Gpt�l t�wh��uj ��S  Y����%  �j�  Y�e� �wh�u�;5��t6��tV�p��u��p�tV�D���Y����Gh�5���u�V�p�E������   뎋u�j�U  YË�U���S3�S�M��F��������u��   ��p8]�tE�M��ap��<���u��   ��p�ۃ��u�E��@��   ��8]�t�E��`p���[�Ë�U��� �p�3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�����   �E��0=�   r����  �p  ����  �d  ��P��p���R  �E�PW�tp���3  h  �CVP�_���3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�����M��k�0�u������u��*�F��t(�>����E�����D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C����Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95��X�������M�_^3�[�{�����jh���"  �M���������}�������_h�u�u����E;C�W  h   �j���Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�p��u�Fh=p�tP� ���Y�^hS�=p���Fp��   �����   j�  Y�e� �C���C���C��3��E��}f�LCf�E�@��3��E�=  }�L����@��3��E�=   }��  ����@���5���p��u���=p�tP�g���Y���S���E������   �0j�  Y��%���u ��p�tS�1���Y�   �    ��e� �E��q!  Ã=, uj��V���Y�,   3�Ë�U��3�9Ev�M�9 t@A;Er�]Ë�U��E3�;͈�tA��-r�H��wjX]Ë͌�]�D���jY;��#���]�������u���Ã���������u���Ã�Ë�U��V������MQ�����Y�������0^]��������������Q�L$+ȃ����Y�z�  Q�L$+ȃ����Y�d�  U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh���:  �e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E��<  Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[��������*3�Ë�U���V�u�M�觘���u�P��  ��e�F�P������Yu��P���  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M��4����E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�0�  �M��E��M��H��EP迸  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�#���@PV�V������^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M�������3�;�u+����j_VVVVV�8�������}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�����j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h�SV�٘����3ۅ�tSSSSS�������N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F�0t�90uj�APQ蕟�����}� t�E��`p�3�_^[�Ë�U���,�p�3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�׸  3ۃ�;�u�y���SSSSS�0脧�������o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q��  ��;�t���u�E�SP�u��V�u��������M�_^3�[�L����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   腔��9}}�}�u;�u+����j^WWWWW�0藦�����}� t�E�`p����  9}vЋE��� 9Ew	�Q���j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�ղ  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� 蝷  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �I�  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�A�����u�E�8 u���} �4����$�p���WF�ն  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP谵  0�F�U�����;�u��|��drj jdRP芵  0��U�F����;�u��|��
rj j
RP�d�  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N������u-�.���j^�03�PPPPP�4������}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V�{������}� t�E��`p�3�_^[�Ë�U���,�p�3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�}�  3ۃ�;�u����SSSSS�0�*��������Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P覱  ��;�t���u�E�SV�u���`������M�_^3�[�����Ë�U���0�p�3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�²  3ۃ�;�u�d���SSSSS�8�o��������   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW��  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[�����Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3��� ��6������Y���(r�_^Ë�Vh   h   3�V趲  ����tVVVVV覞����^Ë�U�������]�����]��E��u��M��m��]����]�����z3�@��3���h���p��th �P�|p��tj ���������U���(3�S�]V�uW�}�E��E��E��E��E��E��E��E�9t�5�*�B���Y��o��M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E����M��]�Q��]���]���Y����  �w���� "   �  �E�����M��]�Q��E�   �]���]���Y�j  �E�   �E�����E�؇��]���]���"  �M��E�؇�r����E�ԇ�׉M��E�ԇ�Z����E��놃�tNIt?It0It ��t����   �E�̇��E�ć��E������E���x����E�   ��������   �E�   �Eܼ���������������   �$��C�E�ԇ��E�؇��E�����Eܴ���Eܬ���Eܤ��y����Eܜ��m����Eܘ���Eܔ���Eܐ���M����]���]�M��]�Q�E�   ��Y��u������ !   �E��_^[���B�BCCCC�B+C�B�B7C@CIC�%�* �G�����*3�Ë�U��QQSV���  V�5(��A�  �EYY�M�ظ�  #�QQ�$f;�uU��  YY��~-��~��u#�ESQQ�$j�i�  ���rVS���  �EYY�d�ES�hs���\$�E�$jj�?�R�  �]��EY�]�Y����DzVS賷  �E�YY�"�� u��E�S���\$�E�$jj�J�  ��^[�Ë�U��QQSV���  V�5,��l�  �EYY�M�ظ�  #�QQ�$f;�uU��  YY��~-��~��u#�ESQQ�$j蔴  ���rVS� �  �EYY�d�ES�hs���\$�E�$jj�?�}�  �]��EY�]�Y����DzVS�޶  �E�YY�"�� u��E�S���\$�E�$jj�u�  ��^[��U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]Ã%�* Ë�U��3�9Ej ��h   P��p���u]�3�@�|*]Ã=|*uWS3�9d*W�=Pp~3V�5h*��h �  j �v���p�6j �5�׃�C;d*|�^�5h*j �5��_[�5��p�% Ë�VW3���<�<�u��8��8h�  �0���p�  YY��tF��$|�3�@_^Ã$�8� 3����S�$pV�8�W�>��t�~tW��W�����& Y����X |ܾ8�_���t	�~uP�Ӄ���X |�^[Ë�U��E�4�8��,p]�jh��  3�G�}�3�9u�TE  j�C  h�   �=:  YY�u�4�8�9t���nj�T���Y��;�u�����    3��Qj
�Y   Y�]�9u,h�  W�g�  YY��uW����Y�����    �]���>�W����Y�E������	   �E��H  �j
�(���YË�U��EV�4�8��> uP�"���Y��uj�19  Y�6�(p^]Ë�U��d*�h*k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �`����   �x*�5�ph @  ��H� �  SQ�֋x*�`�   ���	P�`�@�x*����    �`�@�HC�`�H�yC u	�`��`�x�ueSj �p�֡`�pj �5�Pp�d*�`k��h*+ȍL�Q�HQP�͋���E���d*;`v�m�h*�p*�E�`�=x*[_^�át*V�5d*W3�;�u4��k�P�5h*W�5��p;�u3��x�t*�5d*�h*k�5h*h�A  j�5�`p�F;�t�jh    h   W��p�F;�u�vW�5�Pp뛃N��>�~�d*�F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W��p��u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U����d*�Mk�h*������M���SI�� VW}�����M���������3���U��p*����S�;#U�#��u
���];�r�;�u�h*��S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1�h*�	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t�p*�C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;`u�M�;x*u�%` �M���B_^[����hpTd�5    �D$�l$�l$+�SVW�p�1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q���������������̋�U���S�]V�s35p�W��E� �E�   �{���t�N�38�y���N�F�38�y���E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���@�  �E���|@G�E��؃��u΀}� t$����t�N�38�x���N�V�3:�x���E�_^[��]��E�    �ɋM�9csm�u)�=T� t hT�賨  ����t�UjR�T����M��  �E9Xthp�W�Ӌ���  �E�M��H����t�N�38��w���N�V�3:��w���E��H���y�  �����9S�R���hp�W��葕  �����X á`*Vj^��u�   �;�}�ƣ`*jP�	���YY�@��ujV�5`*����YY�@��ujX^�3ҹX ��@��� �����|�j�^3ҹh W������@����������t;�t��u�1�� B��� |�_3�^������=� t��  �5@�"���YË�U��V�u�X ;�r"���w��+�����Q�����N �  Y�
�� V�(p^]Ë�U��E��}��P������E�H �  Y]ËE�� P�(p]Ë�U��E�X ;�r=�w�`���+�����P�����Y]Ã� P�,p]Ë�U��M���E}�`�����Q����Y]Ã� P�,p]Ë�U��V�uW3�;�u����WWWWW�    蛈������   �F����   �@��   �t�� �F��   ���F�  u	V�  Y��F��v�vV�W  YP��  ���F;���   �����   �F�uOV�-  Y���t.V�!  Y���t"V�  ��V�<�@�  ��Y��Y����@$�<�u�N    �~   u�F�t�   u�F   ��N�A���������	F�~���_^]�jTh8�� ���3��}��E�P��p�E�����j@j ^V�)���YY;��  �@�54��   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@�@��   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j 蛥��YY��tV�M���@��4 ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=4|���=4�e� ��~m�E����tV���tQ��tK�uQ��p��t<�u���������4�@�E� ���Fh�  �FP�ܢ  YY����   �F�E�C�E�9}�|�3ۋ���5@����t���t�N��r�F���uj�X�
��H������P��p�����tC��t?W��p��t4�>%�   ��u�N@�	��u�Nh�  �FP�F�  YY��t7�F�
�N@�����C���g����54��p3��3�@Ëe��E������������Ë�VW�@�>��t1��   �� t
�GP�$p���@   ;�r��6臅���& Y����@|�_^Ë�U��EV3�;�u�����VVVVV�    �τ���������@^]Ë�U��QV�uV�����E�FY��u����� 	   �N ����/  �@t�o���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,������� ;�t�������@;�u�u萫  Y��uV��   Y�F  W��   �F�>�H��N+�I;��N~WP�u�  ���E��M�� �F����y�M���t���t�����������@����@ tjSSQ��  #����t%�F�M��3�GW�EP�u�  ���E�9}�t	�N �����E%�   _[^�Ë�U���dh   �ġ��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U���  �ԏ  �p�3ŉE��EV3���4�����8�����0���9uu3���  ;�u'������0����VVVVV�    跂��������  SW�}�����4�@�����ǊX$�����(�����'�����t��u0�M����u&�a���3��0�E���VVVVV�    �L������C  �@ tjj j �u���  ���u荩  Y����  ��D���  �w����@l3�9H�������P��4�� �����p���`  3�9� ���t���P  ��p��4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P辌  Y��t:��4���+�M3�@;���  j��@���SP�֪  �������  C��D����jS��@���P貪  �������  3�PPj�M�Qj��@���QP�����C��D����hp�����\  j ��<���PV�E�P��(���� �4��p���)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4��p����  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@���迧  Yf;�@����h  ��8����� ��� t)jXP��@���蒧  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4��p���B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4��p���b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �hp��;���   j ��,���P��+�P��5����P��(���� �4��p��t�,���;����Lp��@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0��p��t��,�����@��� ��8�����Lp��@�����8��� ul��@��� t-j^9�@���u�8���� 	   �@����0�?��@����D���Y�1��(�����D@t��4����8u3��$������    � ����  ������8���+�0���_[�M�3�^�.i����jhX��l����E���u������  ����� 	   ����   3�;�|;4r!�����8����� 	   WWWWW�{�����ɋ�����@��������L1��t�P蝦  Y�}���D0t�u�u�u�.������E������� 	   �&����8�M���E������	   �E��������u��  Y�jhx������E���u������ 	   ����   3�;�|;4r����� 	   SSSSS�z�����Ћ����<�@��������L��t�P�Х  Y�]���Dt1�u�D�  YP��p��u�Lp�E���]�9]�t�S����M��6���� 	   �M���E������	   �E�������u��  YË�U��V�u�F��t�t�v�z���f����3�Y��F�F^]Ë�U��   賆  �p�3ŉE�SV�uWV�������3�9FY������}�FjPPS� �  ������������������|��s
������  ������@��������� ��ÊH$����F  ������u�F�������+�ʋǋ��  ��V��+��V���������Z  �������  3�9P0�  �����9Vu�������������<  R�p,�p(�������/�  ��������� Ã���;p(�0���;x,�'���j ������Qh   ������Q�0��p������j �������������������Ξ  ����������������������������;��������������t7������K;�s+���u�J�;�s�H�9
u���������@��uЍ�����+�3����L  �@�t�V��:
u������B;�r������������u�������  ��x������    �$����F��   �V��u!�������   +N��@�����   jj j �������˝  ��;�����u$;�����u�F�8��8
uG@;�r��F    �Yj ������������������胝  �����������������   ;�w�N��t
����   t�~������� �DtG������u��)����������� ������uѭ����������3������������M�_^3�[��c����jh���2����u�����Y�e� �u����Y�E��U��E������   �E��U��D�����u�4���YË�U��V�uV��  Y���u�,���� 	   ����MW�uj �uP��p�����u�Lp�3���tP����Y����������@�����D0� ���_^]�jh���s����E���u������  ����� 	   ����   3�;�|;4r!�����8����� 	   WWWWW�u�����ɋ�����@��������L1��t�P褠  Y�}���D0t�u�u�u��������E���%���� 	   �-����8�M���E������	   �E��������u��  YË�U���SW�}3�;�u �����SSSSS�    ��t��������f  W�����9_Y�E�}�_jSP�������;ÉE�|ӋW��  u+G�.  ��OV��+�u���tA�U��u�����@�����D2�t��;�s���:
u�E�3�B;�r�9]�u�E���   ��x��.����    �   �G��   �W;�u�]��   �]��u�+��������@�E����D0�tyjj �u�������;E�u �G�M��	�8
u�E@;�r��G    �@j �u��u����������}����:�   9Ew�O��t��   t�G�E��D0t�E�E)E��E�M��^_[�Ë�U��V�u�FW��ty�}��t
��t��uh���F��uV�I���EYU3�V�w���FY��y����F��t�t�   u�F   W�u�uV����YP�B�  #����t3��������    ���_^]�jh���^����u�!���Y�e� �u�u�u�u�:������E��E������	   �E��k�����u�[���YË�U��V�uWV�=�  Y���tP�@��u	���   u��u�@Dtj��  j���	�  YY;�tV���  YP� p��u
�Lp���3�V�Y�  ������@����Y�D0 ��tW����Y����3�_^]�jh���s����E���u������  ����� 	   ����   3�;�|;4r!�����8����� 	   WWWWW�q�����ɋ�����@��������L1��t�P褜  Y�}���D0t�u�����Y�E���-���� 	   �M���E������	   �E�������u���  YË�U��9EuF�jP;Mu+�����YY���u3�]ËE�    �6�u�7�e�����Q�/�������tՉ�&3�@]Ë�U���EP�������EYu��߃�]��Jx	�
�A�
�R�����YË�U��}�t]�s��]Ë�U��S�U�������؃��t��P車��Y��u��[]Ë�U����  �p�3ŉE��M�EV3�W�}�������|�����d�����T���ǅ$���^  ��0����������x���;�u �����VVVVV�    ��o��������5  ;�t��@@SuzP�����Y�����t���t�ȃ��������@����A$u&���t���t�ȃ������@����@$�t �V���VVVVV�    �]o��������  �u������]���ƅc��� ��t�����<������k  ��d�����P�x���Y��t0��t���VV��t�������YP�k���YYG�P�M���Y��u��  �<%�1  8G�  3���@���ƅ/��� ��X�����L�����l���ƅa��� ƅ`��� ƅj��� ƅS��� ƅb��� ƅs��� ƅk�����(���G���P�Ƈ��Y��t��l�����L���k�
�DЉ�l�����   ��N��   ��   ��*tp��F��   ��It��Lut��k����   �O��6u�G�84u��(�������4�����8����m��3u�G�82u���\��dtW��itR��otM��xtH��Xu�A��j����9��ht(��lt��wt��S����"�G�8lt���k�����s������k�����s�����S��� �������j��� ��H���u������0�������������3�2ۉ�D���8�s���u�<Stƅs����<Cuƅs������ ��\�����ntJ��ct��{t��d�����t����}���Y���d�����t����@�����x��������  ��D�����H�����L�����t��l��� ��  ��\�����o�r  �  ��c�
  jdZ;���  �z  ��g~E��it!��n�g  ��j��� ��t����f
  �
  ��\�����x���-�4  ƅ`����1  3ۃ�x���-u��T���� -C�	��x���+u��l�����d�����t����^�����x�����L��� u��l������x����k��l�����l�����tf��x�����T�����X������0���P��|���PCS��T�����$�������������
  ��d�����t����������x�����P�̈́��Y��u���������   � � ��a���:�x�����   ��l�����l�������   ��d�����t���������T�����x�����a������0���P��|���PCS��T�����$��������������	  ��x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$����{���������	  ��d�����t����������x�����P�ƃ��Y��u���X��� �_  ��x���et��x���E�I  ��l�����l������5  ��T����e��0���P��|���PCS��T�����$��������������  ��d�����t����D�����x�����-u,��T����-��0���P��|���PCS����������  �	��x���+u/��l�����l�����u!�l������d�����t����������x�����x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$������������  ��d�����t����j�����x�����P�Z���Y��u���d�����t�����x����U�����X��� YY��  ��j��� ��  ��T�����<��������QP��D���� ��k���HP�5�趫��Y�Ѓ��  ��u��l���ǅL���   ��s��� ~ƅb�����d�����t���W��x�����@�������YY��L��� t��l�����l������3  ��t������x�����x�������  ��\���ctN��\���su��	|	����  �� u2��\���{��  ��a���3ҋȃ�B������L�3˅���  ��j��� ��  ��b��� �~  �� �����P��r  Y��t��t������������!��������P�����ǅ���?   ���   �� ���P�����P�֏  f�������f�FF�  ��p��  �������HH�{  ���������t3�;�x�����  ��c�����j��� �  �����������  ��s��� ~ƅb���G�?^��u
�wƅa����j �E�j P�W�����>]u	�]F�E� �f��/����^F<-uB��t>���]t7F:�s�����:�w"*������Ћσ��ǳ�����D�GJu�2���ȊЋ��������D��<]u����  ��H�����D���������x���+u'��l���u��t����d�����t����C�����x���j0^9�x����x  ��d�����t���������x���<xtX<XtT��\���xǅX���   t"��L��� t
��l���u��ǅ\���o   �$  ��d�����t���P�����YY��x����  ��d�����t���������L��� ��x���t��l�����l���}��ǅ\���x   ��   �F��D����������@���������t���WP�j���YY9�@�����  ��j��� �  ��<�����\���c��  ��b��� t��D���3�f���  ��D����  ��  ƅk�����x���-u	ƅ`����	��x���+u'��l���u��t����d�����t���������x�����(��� �J  ���  ��\���xte��\���pt\��x���P�}��Y����   ��\���ou"��x���8��   ��4�����8��������Rj j
��8�����4���茑  �����7��x���P�}��Y��tr��4�����8�����x������������Y��x�����x�����X�����Й����L��� ��4�����8���t��l���t5��d�����t���������x���������d�����t�����x�������YY��`��� ��@�����   ��4�����8����؃� �ى�4�����8�����   ��@�������   ��\���xt;��\���pt2��x���P�1|��Y����   ��\���ou��x���8}n���,k�
�'��x���P�|��Y��tR��x����������Y��x�����X�����L��� ��x����|�t��l���t5��d�����t���������x����X�����d�����t�����x�������YY��`��� t�߃�\���Fu��X��� ��X��� �  ��j��� u8��<�����D�����(��� t��4������8����F���k��� t�>�f�>��H�����c���G��H����`<%u
�G�8%u����t�������������G��x�����H���;�ul��P��l  Y��t!��t�����������G��H���;�uG��t�����x����u�?%uD��H����xnu8������	����*��d�����x�������YY�VS��VP����VS�y�������0���u��T����ra��Y��x����u*��<�����u8�c���u�������� t%������ap������� t
������`p���<���[�M�_3�^��M���Ë�U���VW�u�M��JN���E�u3�;�t�0;�u,�Q���WWWWW�    �X`�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�2  �M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&谱���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9�uh���P������]Ë�U��W��  W�p�u�xp���  ��`�  w��t�_]Ë�U���P  �u�	  �5����h�   �Ѓ�]Ë�U��h���xp��th�P�|p��t�u��]Ë�U���u�����Y�u��p�j�5���Y�j�R���YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=(| th(|��z  Y��t
�u�(|Y�
���h�qhxq����YY��uBhډ��o���\q�$tq�c����=0 Yth0�z  Y��tj jj �03�]�jh��Q���j�Q���Y�e� 3�C9���   ���E���} ��   �5(蝟��Y���}؅�tx�5$舟��Y���u܉}�u����u�;�rW�d���9t�;�rJ�6�^������N�������5(�H������5$�;�����9}�u9E�t�}�}؉E����u܋}��h�q��q�_���Yh�q��q�O���Y�E������   �} u(��j����Y�u�����3�C�} tj�f���Y��w���Ë�U��j j�u�������]�jj j ������Ë�V腞����V��  V�x  V�"Z��V��  V�щ  V�3  V�L��V�p���hׄ�ם����$�^Ã=, u腭��V�5lW3���u����   <=tGV�z��Y�t���u�jGW�y����YY�=x��tˋ5lS�BV�vz����C�>=Yt1jS�wy��YY���tNVSP�'K������t3�PPPPP�kY�������> u��5l��Z���%l �' �    3�Y[_^��5x��Z���%x ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�Ո  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#���  Y��t��M�E�F��M��E���͇  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9,u����h  ��VS����p��*�5�;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�v����Y;�t)�U��E�P�WV�}�������E���H�l�5p3�����_^[�Ë�U�졨��SV�5�pW3�3�;�u.�֋�;�t��   �#�Lp��xu
jX���������   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5hpSSS+�S��@PWSS�E��։E�;�t/P��u��Y�E�;�t!SS�u�P�u�WSS�օ�u�u��W��Y�]��]�W��p���\��t;�u���p��;��r���8t
@8u�@8u�+�@P�E��gu����Y;�uV��p�E����u�VW�K����V��p��_^[�Ë�V�,��,�W��;�s���t�Ѓ�;�r�_^Ë�V�4��4�W��;�s���t�Ѓ�;�r�_^Ë�U��QQV�X��������F  �V\�(W�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ��= ���;�}$k��~\�d9 �=� B߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]Ë�U����p��e� �e� SW�N�@��  ��;�t��t	�Уt��`V�E�P�q�u�3u�� q3��Xp3���p3��E�P��p�E�3E�3�;�u�O�@����u������5p��։5t�^_[�Ë�U��QQS�]VW3�3��}�;�0t	G�}���r���w  j茄  Y���4  j�{�  Y��u�=x�  ���   �A  h0��  S��W�aD������tVVVVV�R����h  ��Vj �� ��p��u&h�h�  V�D������t3�PPPPP�cR����V�1s��@Y��<v8V�$s����;�j��h�+�QP� :  ����t3�VVVVV� R�����3�h�SW�69  ����tVVVVV��Q�����E��4�4SW�9  ����tVVVVV��Q����h  h�W��  ���2j���p��;�t$���tj �E�P�4�4�6�or��YP�6S��p_^[��j��  Y��tj��  Y��u�=xuh�   �)���h�   ����YYË�U��E��]Ë�U���5��y���Y��t�u��Y��t3�@]�3�]��A@t�y t$�Ix��������QP�Y���YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u蛤���8*u�ϰ?�d����} �^[]Ë�U���x  �p�3ŉE�S�]V�u3�W�}�u��������������������������������������������������������������>����u5�����    3�PPPPP�Q���������� t
�������`p������
  �F@u^V�����Y�����t���t�ȃ��������@����A$u����t���t�ȃ������@����@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw����H���3��3�3����h�j��Y������;���	  �$�O���������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�������/Y  Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u��������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P�~  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  ��������P�~k��Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7���������|  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V�?i��������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5��m���Y�Ћ���������   t 9�����u������PS�5$��>���Y��YY������gu;�u������PS�5 �����Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�v  ��0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u���������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF�/y  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t��������F�������� Y���������������t������������������������� t
�������`p��������M�_^3�[�p3���ÐZ�[����5�@�������U���   �p�3ŉE��ESV�u3ۃ}W��t�����l�����   Sh�   ��|�����Q�u��x����uP�oy  ����;�uj�Lp��z��   SSS�u�u��t����Cy  ����p���;�t_3�FVP�)d����YY;�tMS��p�����x���W�u�u��t����y  ����;�tjV��c��YY��l����;�u!9�x���tW�E��Y����M�_^3�[�N2���ÍN�QWVP�+  ����tSSSSS�C����9�x���tW�UE��Y3��9]u�Sj��W�u�uP�w  ����t�����P��]��Y��tɊ�
���,0GG����|�뱋�U��E��]�jh8������3��]3�;���;�u�<����    WWWWW�CD��������S�=|*u8j�ɬ��Y�}�S����Y�E�;�t�s���	�u���u��E������%   9}�uSW�5�q����迷���3��]�u�j藫��Y�U���0���S�ٽ\�����=� t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=� t�#  ��8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����,  �   [�À�8�����=\ uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �������������؎����s4����,ǅr���   ��������������Ў����v���VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P��u  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����D   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Àzuf��\���������?�f�?f��^���٭^�����剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-���p��� ƅp���
��
�t����������l$�l$�D$���   5   �   t�������  u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t�0���0���l$����4���4���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r �������8�|$�l$�ɛ�l$������l$��Ã�,��?�$�~����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  ������< �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����l�Ƀ�u�\$0�|$(���l$�-t�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�\�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���T�|$�T�<$� �|$$�D$$   �D$(�l$(���T�<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  ������< �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����l�Ƀ�u�\$0�|$(���l$�-t�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�\�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���T�|$�T�<$� �|$$�D$$   �D$(�l$(���T�<$�l$$�Q�����0Z�����0Z�������@���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�e  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   �� ��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��,������������������   s��<���$������������������   v��4�떋�U����p�3ŉE�j�E�Ph  �u�E� �q��u����
�E�P�E=��Y�M�3��	���Ë�U���4�p�3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5tp�M�QP�֋lp��t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u���N����YF;�~[�����wS�D6=   w/�T�����;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�?��Y;�t	� ��  ���E���}�9}�t؍6PW�u������V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�hp��t`�]��[�hp9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�M��YY�E�;�t+WWVPV�u�W�u��;�u�u��.��Y�}���}��t�MЉ�u�����Y�E��e�_^[�M�3��U���Ë�U���S�u�M�����]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P��8  YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP��  �� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U��QQ�p�3ŉE���SV3�W��;�u:�E�P3�FVh(}V�q��t�5��4�Lp��xu
jX���������   ;���   ����   �]�9]u��@�E�5lp3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w������;�t� ��  �P�<��Y;�t	� ��  ���؅�ti�?Pj S�?����WS�u�uj�u�օ�t�uPS�u�q�E�S�����E�Y�u3�9]u��@�E9]u��@�E�u�����Y���u3��G;EtSS�MQ�uP�u��������;�t܉u�u�u�u�u�u�q��;�tV�-,��Y�Ǎe�_^[�M�3������Ë�U����u�M��N���u$�M��u �u�u�u�u�u�������}� t�M��ap���jhX��ߞ���M3�;�v.j�X3���;E�@u�~���    WWWWW�+����3���   �M��u;�u3�F3ۉ]���wi�=|*uK������u�E;l*w7j�q���Y�}��u�w���Y�E��E������_   �]�;�t�uWS�����;�uaVj�5�`p��;�uL9=�t3V����Y���r����E;��P����    �E���3��uj����Y�;�u�E;�t�    �������jhx�������]��u�u�J:��Y��  �u��uS�*��Y�  �=|*��  3��}�����  j�~���Y�}�S角��Y�E�;���   ;5l*wIVSP艗������t�]��5V�X���Y�E�;�t'�C�H;�r��PS�u�����S�W����E�SP�}�����9}�uH;�u3�F�u������uVW�5�`p�E�;�t �C�H;�r��PS�u��w��S�u��0������E������.   �}� u1��uF������uVSj �5��p����u�]j诐��YË}����   9=�t,V�h���Y��������{��9}�ul���LpP�V{��Y��_����   �{��9}�th�    �q��uFVSj �5��p����uV9�t4V�����Y��t���v�V�����Y�:{���    3�� �����'{���|�����u�{�����LpP��z���Y���ҋ�U��MS3�;�v(j�3�X��;Es��z��SSSSS�    ��'����3��A�MVW��9]t�u�[���Y��V�u������YY��t;�s+�Vj �S�������_^[]Ë�U��E��������]Ë�U��E�(V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5��aj��Y�j h���ɚ��3��}�}؋]��Lt��jY+�t"+�t+�td+�uD��k�����}؅�u����a  �����`�w\���]���������Z�Ã�t<��t+Ht�y���    3�PPPPP�&����뮾���������
�����E�   P�i���E�Y3��}���   9E�uj�����9E�tP����Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.��M܋ ��9M�}�M�k��W\�D�E����i����E������   ��u�wdS�U�Y��]�}؃}� tj 聍��Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3��k���Ë�U����HB�PD�M��U���u����Ãe� SW�E��FPj1Q3�C�E�SP�P������FPj2�u��E�SP�;�����FPj3�u��E�SP�&�����FPj4�u��E�SP������P��FPj5�u��E�SP�������FPj6�u��E�SP�����Vj7�u���E�SP�������F Pj*�u��E�SP������P��F$Pj+�u��E�SP������F(Pj,�u��E�SP������F,Pj-�u��E�SP�{�����F0Pj.�u��E�SP�f�����P��F4Pj/�u��E�SP�N�����FPj0�u��E�SP�9�����F8PjD�u��E�SP�$�����F<PjE�u��E�SP������P��F@PjF�u��E�SP�������FDPjG�u��E�SP�������FHPjH�u��E�SP�������FLPjI�u��E�SP������P��FPPjJ�u��E�SP������FTPjK�u��E�SP������FXPjL�u��E�SP�v�����F\PjM�u��E�SP�a�����P��F`PjN�u��E�SP�I�����FdPjO�u��E�SP�4�����FhPj8�u��E�SP������FlPj9�u��E�SP�
�����P��FpPj:�u��E�SP�������FtPj;�u��E�SP�������FxPj<�u��E�SP�������F|Pj=�u��E�SP������P����   Pj>�u��E�SP��������   Pj?�u��E�SP��������   Pj@�u�S�E�P�h�������   PjA�u��E�SP�P�����P����   PjB�u��E�SP�5�������   PjC�u��E�SP��������   Pj(�u��E�SP��������   Pj)�u��E�SP�������P����   Pj�u��E�SP���������   Pj �u��E�SP��������   Ph  �u��E�SP��������   Ph	  �]�S�E�j P������P���_���   [�Ë�U��V�u����  �v��!���v��!���v��!���v��!���v�!���v�!���6�!���v �!���v$�!���v(�!���v,�!���v0�!���v4�}!���v�u!���v8�m!���v<�e!����@�v@�Z!���vD�R!���vH�J!���vL�B!���vP�:!���vT�2!���vX�*!���v\�"!���v`�!���vd�!���vh�
!���vl�!���vp�� ���vt�� ���vx�� ���v|�� ����@���   �� �����   �� �����   � �����   � �����   � �����   � �����   � �����   � �����   �| �����   �q �����   �f ����,^]Ë�U��SVW�}�  ��t@h�   j�}>����YY��u3�@�E��������tV�+���V� ��YY��ǆ�      �����   �;�t�   P�p�73�_^[]Ë�U��V�u��t5�;@tP����Y�F;DtP���Y�v;5HtV���Y^]Ë�U���S�]V3�W�]�u�9su9su�u��u��E@�:  j0j�=����YY�};�u3�@�w  ���   jYj��<=��3�Y�E�;�u�u�0��Y�щ09s��   j�=��Y�E�;�u3�F�u����u�� ��YY���  �0�u�{>VjW�E�jP�[����E�FPjW�E�jP�F���	E�FPjW�E��E�jP�.�����<E�tV����Y���뎋E�� ����0|��9��0�@�8 u��7��;u���~�����> u���@�E��D�H�H�u��H�E�3�A��E���t����   �5p��tP�֋��   ��tP�օ�u���   ������   ����YY�E����   �E����   �E���   3�_^[�Ë�U��V�u��t~�F;LtP���Y�F;PtP���Y�F;TtP���Y�F;XtP���Y�F;\tP�r��Y�F ;`tP�`��Y�v$;5dtV�N��Y^]Ë�U���SV�uW3��}��u��}�9~u9~u�}��}��@�6  j0j�M;����YY;�u3�@�u  j��:��Y�E�;�u	S����Y���89~��  j��:��Y�E�;�uS�����u����Y�҉8�v8�CPjV�E�jP�������CPjV�E�jP������CPjV�E�jP�������CPjV�E�jP�������P��CPjV�E�jP�������C PjPV�E�jP������C$PjQV�E�jP������C(PjV�E�j P������P��C)PjVj �E�P�y�����C*PjTV�E�j P�e�����C+PjUV�E�j P�Q�����C,PjVV�E�j P�=�����P��C-PjWV�E�j P�&�����C.PjRV�E�j P������C/PjSV�E�j P�������<�t$S����S�o���u��g���u��_�����Q����C����0|��9��0�@�8 u��#��;u���~�����> u���jY�@���E�u�   ��	���I�K� �@�M��C3�@3��9}�t�M�����   ;�tP�p���   ;�t#P�p��u���   ������   ���YY�E����   �E����   ���   3�_^[��3�Ë�U��ES3�VW;�t�};�w��l��j^�0SSSSS���������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u��l��j"Y����3�_^[]�����������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^�Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w��k��j^�0SSSSS����������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x�����xk��j"Y���낋�U��3�S3�@9]|FVW��t>�EÙ+��E���<��7�E�0�N  YY��u
�M���9�}N�u��^;]~�_^3Ʌ���[��]Ë�U����p�3ŉE�V���tS�> tNhT�V�c��YY��t=hP�V�	c��YY��uj�E�Pj�w�q��t/�u�V�B%��Y�M�3�^�����j�E�Ph  �w�q��u3��׍E�hL�P�b��YY��u���p뻋�U��3�f�Mf;�8�t@@��r�3�@]�3�]Ë�V3��#��,aB<w������,A<w��������tЊ
��u׋�^�3��
B��A|��Z~��a��w@��Ë�U���|�p�3ŉE�VW�}�^\�����ׁƜ   ������jx�E�P�F���%���  PW�q��u!F@�2�E�P�v��L  YY��uW����Y��t
�N�~�~�F���Ѓ��M�_3�^������ ��U���|�p�3ŉE�Vjx�E�P�E%�  j   P���q��u3��.�U������9Et�} t�6W�������V����5��Y;�_t�3�@�M�3�^�N���Ë�U���|�p�3ŉE�SVW�}�Q[�����ׁƜ   �y����q��jx�E�P�F���%���  PW�Ӆ�u�f 3�@�b  �E�P�v��K  YY����   jx�E�P�F���%���  PW�Ӆ�t��E�P�6�K  YY��u�N  �~�R�FuO�F��t,P�E�P�6��L  ����u�6�N�~��4��Y;Fu!�~��V��uW����Y��t	���V�~�N�   #�;���   jx�E�P�F���%���  PW�Ӆ������E�P�6�	K  Y3�Y��u/�N   �F9^t
   �F�G9^t;�6�=4��Y;Fu.j�9^u49^t/�E�P�6�J  YY��uSW�������YY��t�N   9^u�~�F���Ѓ��M�_^3�[�~���� ��U���|�p�3ŉE�VW�}�Y�����ׁƜ   ������jx�E�P�F���%���  PW�q��u!F@�[�E�P�6�J  YY��u	9Fu0j��~ u0�~ t*�E�P�6��I  YY��uPW���$���YY��t
�N�~�~�F���Ѓ��M�_3�^� ���� �6�3���v�����@�F�3��������f @�~ YY�FtjX���	���jhp��F�q�F�   t�   t�u�f ��6�2�������@Y�FtjX������jhB��F�q�Fu�f Ë�U��SVW�+X���]���Ɯ   ��u�N  �   �C@�~����t�8 tWjh�����������f ��tS�8 tN���t�8 t�������S����~ ��   Vj@hx���������tb�?��t�? t�����P�����I�?��t0�? t+W��1������Y�j@hd��F�q�Fu�f ��F  �q�F�F�~ ��   �˃����#ˋ��������}����   ����  ��   ����  ��   ��P��p����   j�v� q����   �E��tf�Nf�f�Nf�Hf�x�]��tm�=q�  f9u%hX�j@S�������t"3�PPPPP�������j@Sh  �v�ׅ�t,j@�C@Ph  �v�ׅ�tj
j��S�u�I  ��3�@�3�_^[]Ë�U��VW�}�ǃ� ��  H��  H��  H�I  H��  �M�ESj Z�r  �0;1t|�0�+�t3ۅ��Í\�����i  �p�Y+�t3ۅ��Í\�����H  �p�Y+�t3ۅ��Í\�����'  �p�Y+�t3ۅ��Í\����3����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3����r  �p;qt~�p�Y+�t3ۅ��Í\�����I  �p	�Y	+�t3ۅ��Í\�����(  �p
�Y
+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����w  �p�Y+�t3ۅ��Í\����3����R  �p;qt~�Y�p+�t3ۅ��Í\�����)  �p�Y+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����x  �p�Y+�t3ۅ��Í\�����W  �p�Y+�t3ۅ��Í\����3����2  �p;qt~�p�Y+�t3ۅ��Í\�����	  �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\����3�����   �p;qtr�p�Y+�t3ۅ��Í\����u}�p�Y+�t3ۅ��Í\����u`�p�Y+�t3ۅ��Í\����uC�p�Y+�t3ۅ��Í\����3���u"��+�;�������σ���  �$�������  �P�;Q�tq���Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����3����v����P�;Q�t}���Q�+�t3҅��T�����N����p��Q�+�t3҅��T�����-����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����}����p��Q�+�t3҅��T����3����X����P�;Q�t}���Q�+�t3҅��T�����0����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T�����^����p��Q�+�t3҅��T����3����9����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�to���Q�+�t3҅��T���u6�p��Q�+�t3҅��T���u�p��Q�+�t3҅��T���t����@��I�+�t3Ʌ����L	����3���u3�[�S  �P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����n����p��Q�+�t3҅��T�����M����p��Q�+�t3҅��T�����,����p��Q�+�t3҅��T����3��������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����x����P�;Q�t}���Q�+�t3҅��T�����P����p��Q�+�t3҅��T�����/����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3����Z����P�;Q�t~�Q��p�+�t3҅��T�����1����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����`����p��Q�+�t3҅��T����3����;����I��@�+�� ���3Ʌ����L	���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����b����p��Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����l����P�;Q�t}���Q�+�t3҅��T�����D����p��Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����s����p��Q�+�t3҅��T����3����N����P�;Q�t~�Q��p�+�t3҅��T�����%����Q��p�+�t3҅��T���������Q��p�+�t3҅��T����������Q��p�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T����3����/���f�P�f;Q�������Q��p�+������3҅��T����  �����P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����i����P�;Q�t}���Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����p����p��Q�+�t3҅��T����3����K����P�;Q�t}���Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T�����r����p��Q�+�t3҅��T�����Q����p��Q�+�t3҅��T����3����,����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T�����3����p��Q�+�t3҅��T����3��������p��Q�+������3҅��T���������������M�u��+�t3҅��T�����   �A�V+�t3҅��T�����   �A�V+�t3҅��T�����   �A�N+���   3Ʌ����L	����   �M�u��+�t3҅��T���uh�A�V+�t3҅��T���uK�A�N랋M�u��+�t3҅��T���u �A�N�p����E�M� �	�_���3�_^]�8�*�6�W���������,���9���|�����������~�^�j�����������l�@�L�l����������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U����SV�uW3��E��}�}��}��FFf�> t����at8��rt+��wt�L��WWWWW�    ������3��S  �  �3ۃM��	�	  �M�3�AFF�f;���  � @  ;��   ����S��   ��   �� ��   ��tVHtG��t1��
t!���u���9}���   �E�   ����   �ˀ   �   ��@��   ��@�   �E�   �   ����   �E����������   �E��}9}�ur�E�   �� �l��TtX��tCHt/��t��������� �  uC��E9}�u:�e������E�   �09}�u%	U��E�   ��� �  u�� �  ��   ��t3���FF�f;������9}���   �FFf�> t�jVhl���:  �����`���j ��X�FFf9t�f�>=�G���FFf9t�jht�V��9  ����u��
��   �Djh��V��9  ����u����   �%jh��V�9  �������������   �FFf�> t�f9>�����h�  �u�ES�uP�p8  ����������E�d�M��H�M�x�8�x�x�H_^[��jh����j��3�3��}�j��_��Y�]�3��u�;5`*��   �@��9t[� �@��uH� �  uA�F���w�FP��^��Y����   �@�4�V�m��YY�@���@�tPV��m��YYF둋��}��h��j8�9��Y�@��@�9tIh�  � �� P�W  YY���@u�4����Y�@����� P�(p�@�<�}�_;�t�g �  �_�_��_�O��E������   ���j��Ë}�j��]��Y�SVW�T$�D$�L$URPQQh��d�5    �p�3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�R  �   �C�d  �d�    ��_^[ËL$�A   �   t3�D$�H3������U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�  3�3�3�3�3���U��SVWj j h��Q�]  _^[]�U�l$RQ�t$������]� ��U����u�M������E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U��3�@�} u3�]�U��SVWUj j h��u�]  ]_^[��]ËL$�A   �   t2�D$�H�3�����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�d�5    �p�3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�u�Q�R9Qu�   �SQ���SQ���L$�K�C�kUQPXY]Y[� ����������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �������U��W�}3�������ك��E���8t3�����_�Ë�U���SV�u�M������]�   ;�sT�M胹�   ~�E�PjS�����M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�h���YY��t�Ej�E��]��E� Y��E��� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�	����$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=� u�E�H���w�� ]�j �u�����YY]Ë�U���(�p�3ŉE�SV�uW�u�}�M��8����E�P3�SSSSW�E�P�E�P�1?  �E�E�VP�4  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�8����Ë�U���(�p�3ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P�>  �E�E�VP�89  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�����Ë�U��MSV�u3�W�y;�u�C��j^�0SSSSS���������   9]v݋U;ӈ~���3�@9Ew��B��j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�F��@PWV�=�����3�_^[]Ë�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���H���u��P������Ɂ���  �P���t�M�_^f�H[�Ë�U���0�p�3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��UC  �uЉC�E։�EԉC�E�P�uV�������$��t3�PPPPP�&������M�_�s^��3�[������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�!���YË�U��E�M%����#�V������t1W�}3�;�tVV�#L  YY���?��j_VVVVV�8���������_��uP�u��t	��K  ����K  YY3�^]Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u�Hp�M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�}  Y����  �t�Etj�c  Y����v  ����   �E��   j�A  �EY�   #�tT=   t7=   t;�ub��M�������{L�H��M�����{,���2��M�����z�����M�����z�������������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�x  �M��]�� �����������}�E���@{�S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}�:��� "   ]��:��� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3��Ř;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P��������uV�,���Y�E�^�ËŜ�h��  �u(�  �u�����E ���Ë�U��=� u(�u�E���\$���\$�E�$�uj�/�����$]��9��h��  �u� !   �J  �EYY]Ë�S��QQ�����U�k�l$���   �p�3ŉE��s �CP�s��������u"�e���CP�CP�s�C �sP�E�P�I������s�p������=� u+��t'�s �C���\$���\$�C�$�sP�r�����$�P�����$��  �s �  �CYY�M�3�������]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj���  f;�u�E�� u9Utj��3�]Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������"Q���EQQ�$����������  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�-��]���t����-��]�������t
�-��]����t	�������؛�� t���]����jh���MW��3�9�*tV�E@tH9�t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%� �e��U�E�������e��U�-W��Ë�U��E�4]�jh����V���e� �u�u�$q�E��/�E� � �E�3�=  �����Ëe�}�  �uj��p�e� �E������E��V��Ë�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h�hpTd�    P��SVW�p�1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh8��U��3ۉ]�j�J��Y�]�j_�}�;=`*}W�����@�9tD� �@�tP�����Y���t�E��|(�@��� P�$p�@�4����Y�@�G��E������	   �E���T���j�H��YË�U����UV�uj�X�E�U�;�u��3���  �3��� 	   ����  S3�;�|;54r'�3����3��SSSSS� 	   ����������Q  ����W�<�@�����ƊH��u�`3����F3��� 	   �j�����wP�]�;��  ����  9]t7�@$����E���HjYtHu���Шt����U�E�E��   ���Шu!��2�����2���    SSSSS��������4����M;�r�E�u�B���Y�E�;�u�2���    �2���    ����h  jSS�u�^  ��D(�E���T,���AHtt�I��
tl9]tg��@�M�E�   �D
8]�tN��L%��
tC9]t>��@�M�}��E�   �D%
u$��L&��
t9]t��@�M�E�   �D&
S�M�Q�uP��4��p���{  �M�;��p  ;M�g  �M��D� ���  �}��  ;�t�M�9
u��� ��]�E�É]�E�;���   �M�<��   <t�CA�M�   �E�H;�s�A�8
u
AA�M�
�u�E�m�Ej �E�Pj�E�P��4��p��u
�Lp��uE�}� t?��DHt�}�
t����M��L�%;]�u�}�
t�jj�j��u�  ���}�
t�C�E�9E�G������D� @u����C��+E�}��E���   ����   K���xC�   3�@�����;]�rK�@��� t��������u�M0��� *   �zA;�u��@���AHt$C���Q|	���T%C��u	���T&C+���ؙjRP�u��  ���E�+]���P�uS�u�j h��  �lp�E���u4�LpP��/��Y�M���E�;EtP�R���Y�E�����  �E��  �E��3�;�����E��L0��;�t�M�f�9
u��� ��]�E�É]�E�;���   �E�f����   f��tf�CC@@�E�   �M����;�s�Hf�9
u���Ej
�   �M�   �Ej �E�Pj�E�P��4��p��u
�Lp��u[�}� tU��DHt(f�}�
t�jXf���M��L��M��L%��D&
�*;]�uf�}�
t�jj�j��u�|  ��f�}�
tjXf�CC�E�9E�������t�@u��f� f�CC+]�]������Lpj^;�u�F.��� 	   �N.���0�i�����m�Y����]��\���3�_[^��jhX��N���E���u�.���  ��-��� 	   ����   3�;�|;4r!��-���0��-��� 	   VVVVV��������ɋ�����@��������L9��t�����;M�Au�-���0�-���    �P��  Y�u���D8t�u�u�u�~������E���O-��� 	   �W-���0�M���E������	   �E��N����u�  YË�U��QQ�EV�u�E��EWV�E���  ���Y;�u��,��� 	   �ǋ��J�u�M�Q�u�P��p�E�;�u�Lp��t	P��,��Y�ϋ�����@�����D0� ��E��U�_^��jhx��<M������u܉u��E���u�,���  �p,��� 	   �Ƌ���   3�;�|;4r!�a,���8�G,��� 	   WWWWW�N������ȋ�����@��������L1��u&� ,���8�,��� 	   WWWWW������������[P�=  Y�}���D0t�u�u�u�u�������E܉U���+��� 	   ��+���8�M���M���E������   �E܋U��L����u�z  YË�U��E���u�o+��� 	   3�]�V3�;�|;4r�Q+��VVVVV� 	   �X�����3���ȃ�����@���D��@^]Ë�U����p�3ŉE�V3�95�tO�=�	�u�>:  ��	���u���  �pV�M�Qj�MQP�0q��ug�=�u��Lp��xuω5�VVj�E�Pj�EPV�,qP�hp��	���t�V�U�RP�E�PQ�(q��t�f�E�M�3�^���������   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M������E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P�0���YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�lp���E�u�M;��   r 8^t���   8]��e����M��ap��Y����)��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�lp���:���뺋�U��j �u�u�u�������]Ë�U��EVW��|Y;4sQ���������<�@����<�u5�=xS�]u�� tHtHuSj��Sj��Sj��4q��3�[��(��� 	   ��(���  ���_^]Ë�U��MS3�;�VW|[;4sS������<�@�������@t5�8�t0�=xu+�tItIuSj��Sj��Sj��4q���3���5(��� 	   �=(������_^[]Ë�U��E���u�!(���  �(��� 	   ���]�V3�;�|";4s�ȃ�����@����@u$��'���0��'��VVVVV� 	   ������������ ^]�jh���KH���}����������4�@�E�   3�9^u6j
�&=��Y�]�9^uh�  �FP�0���YY��u�]��F�E������0   9]�t����������@�D8P�(p�E��H���3ۋ}j
��;��YË�U��E�ȃ�����@���DP�,p]�jh���G���M��3��}�j�;��Y��u����b  j�g<��Y�}��}؃�@�<  �4�@����   �u���@   ;���   �Fu\�~ u9j
�<��Y3�C�]��~ uh�  �FP�$���YY��u�]���F�e� �(   �}� u�^S�(p�FtS�,p��@낋}؋u�j
��:��YÃ}� u��F��+4�@��������u�}��uyG�+���j@j ����YY�E���ta��@��4 ���   ;�s�@ ���@
�` ��@�E������}�����σ�����@�DW�����Y��u�M���E������	   �E��EF���j�%:��Y��������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U��E�8]Ë�U����u�M��%����E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U���SVW�
���e� �=< ����   h���8q�����*  �5|ph��W�օ��  P�T���$p�W�<��P�?���$\�W�@��P�*���$@�W�D��P���Y�L��th(�W��P����Y�H�H;�tO9LtGP�[���5L���N��YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9�@;�t0P���Y��t%�ЉE���t�D;�tP����Y��t�u��ЉE��5<����Y��t�u�u�u�u����3�_^[�Ë�U��MV3�;�|��~��u�t�(�t�t��P"��VVVVV�    �W��������^]áp���3�9P����Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v��!��j^SSSSS�0����������V�u�M�蠼���E�9X��   f�E��   f;�v6;�t;�vWSV蚿�����!��� *   �!��� 8]�t�M��ap�_^[��;�t2;�w,�a!��j"^SSSSS�0�i�����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�hp;�t9]�^����M;�t����Lp��z�D���;��g���;��_���WSV�þ�����O�����U��j �u�u�u�u�|�����]Ë�U����u�M��g����u�u�u�u�<q�}� t�M��ap��Ë�U��QQ�p�3ŉE��TS�<qVW3�3�G;�u,VVWV�Ӆ�t�=T�/�Lp��xu
jX�T��T����   ;���   ;�u#9uu�E� �@�EVV�u�u�ӋȉM�;�u3��   ~Ej�3�X���r9�D	=   w�	 ����;�t����  ���P�����Y;�t	� ��  �����3�;�t��u�W�u�u�Ӆ�t VV9uuVV��u�uj�WV�u�hp��W����Y����u�u�u�u�q�e�_^[�M�3�艹���Ë�U����u�M�������u�E��u�u�u�uP�������}� t�M��ap��Ë�S��QQ�����U�k�l$���   �p�3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|�����������uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�(�����h��  ��x��������>YYt�=� uV�ް��Y��u�6�����Y�M�_3�^������]��[Ë�U��UV�uW��H�F��w�� �
�y�B��w�� ��t;�t�_+�^]Ë�U���S�u�M��>���3�9]u.�P��SSSSS�    �W�����8]�t�E��`p������   W�};�u+���SSSSS�    �!�����8]�t�E��`p������U�E�9XuW�u�:���YY�4V�E� �M�QP�����E����M�QP�������G;�t;�t�+���^8]�t�M��ap�_[�Ë�U��V3�95�u09uu���VVVVV�    �����������9ut�^]����V�u�u�������^]Ë�U���S3�VW9]��   �u�M��
���9]u.���SSSSS�    �%�����8]�t�E��`p������   �};�t˾���9uv(����SSSSS�    �������8]�t�E��`p����`�E�9Xu�uW�u�N+  ��8]�tD�M��ap��;�E� �M�QP������E����M�QP������G�Mt;�t;�t�+����3�_^[�Ë�U��V3�95�u99uu�=��VVVVV�    �D����������'9ut܁}���w�^]�*  V�u�u�u������^]Ë�U��QSV��3�;�u����j^SSSSS�0����������   W9]w����j^SSSSS�0����������   3�9]���A9Mw	���j"�ЋM�����"w��]���9]t�-�N�E�   �؋�3��u��	v��W���0�A�E�3�;�v�U9U�rڋE�;Er�럈I���I�G;�r�3�_^[�� ��U��}
�Eu
��}jj
�j �u�u�M�����]Ë�U���4S3��E�VW���]��]��E�   �]�t	�]��E��
�E�   �]��E�P�*,  Y��tSSSSS�������M� �  ��u�� @ u9E�t�M������+ú   ��   �tGHt.Ht&�w������Z��j^SSSSS�0�b������  �U����t��   u��E�   @��}��EjY+�t7+�t*+�t+�t��@u�9}����E���E�   ��E�   ��E�   ��]��E�   #¹   ;��   ;t0;�t,;�t=   ��   =   �@����E�   �/�E�   �&�E�   �=   t=   t`;������E�   �E�E�   ��t�h��#M��x�E�   �@t�M�   �M�   �M��   t	}�� t�M�   ��E�   릨t�M�   �%�������u�����������    �   �E�=@qS�u��    �u�E�P�u��u��u�׉E���um�M��   �#�;�u+�Et%�e����S�u�E��u�P�u��u��u�׉E���u4�6������@�����D0� ��LpP���Y�S��� �u  �u���p;�uD�6������@�����D0� ��Lp��V�<��Y�u�� p;�u�����    룃�u�M�@�	��u�M��u��6������Ѓ�����@Y��Y�M����L��Ѓ�����@���D$� ��M��e�H�M���   �����  �Etrj���W�6�0M�����E�;�u�z���8�   tN�6��P�������j�E�P�6�]��e�������uf�}�u�E�RP�6�/&  ��;�t�SS�6��L����;�t��E���0  � @ � @  �}u�E�#�u	M�	E�E#�;�tD=   t)= @ t"=   t)= @ t"=   t= @ u�E���M�  #�;�u	�E���]��E   ��  �E�@�]���  �E��   �#�=   @��   =   �tw;���  �E�;��y  ��v��v0���f  �E�3�H�&  H�R  �E���  �E�   �  jSS�6��������t�SSS�6�����#���������j�E�P�6����������t�����tk����   �}�﻿ uY�E���   �E�;���   ���b������P���jSS�6�l�������C���SSS�6�W�����#����   �����E�%��  =��  u�6��N��Y�G��j^�0���d  =��  uSj�6��J�������������E��ASS�6��J������E�﻿ �E�   �E�+�P�D=�P�6� E������������9}�ۋ������@�����D$�2M���0�������@�����D$�M�������
ʈ8]�u!�Et��ȃ�����@���D� �}��   ���#�;�u|�Etv�u�� pS�u�E�jP�u������W�u�@q���u4�LpP�>����ȃ�����@���D� ��6�P���Y�����6������@�������_^[��jh���t3��3��u�3��};���;�u���j_�8VVVVV趿�������Y��3�9u��;�t�9ut�E%������@tu��u�u�u�u�E�P���i������E��E������   �E�;�t���-3���3��}9u�t(9u�t�����������@�D� ��7�����YË�U��j�u�u�u�u�u������]Ë�U���SV3�3�W9u��   �];�u"����VVVVV�    �ɾ���������   �};�t��u�M��u����E�9pu?�f��Ar	f��Zw�� ���f��Ar	f��Zw�� CCGG�M��tBf��t=f;�t��6�E�P�P��#  ���E�P�P��#  ��CCGG�M��t
f��tf;�t�����+��}� t�M��ap�_^[�Ë�U��V3�W95�u3�9u��   �};�u����VVVVV�    �۽���������`�U;�t��f��Ar	f��Zw�� ���f��Ar	f��Zw�� GGBB�M��t
f;�tf;�t�����+��V�u�u�u�w�����_^]Ë�U��} u3�]ËU�M�Mt�f��tf;uAABB����
+�]Ë�U����  ��f9Eu�e� �e�   f9Es�E��f�Af#E���E��@�u�M�踪���E��p�p�E�Pj�EP�E�jP�#  ����u!E��}� t�E�`p��E��M#��Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�	N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC��	��+�	;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�	N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���	A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�	��	��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}础	��	�3�@�   ��	�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+�	��M���Ɂ�   �ً�	]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�	N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC��	��+�	;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�	N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���	A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;�	��	��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}硘	��	�3�@�   ��	�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+�	��M���Ɂ�   �ً�	]���@u�M�U�Y��
�� u�M�_[�Ë�U���|�p�3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u���SSSSS�    �ı����3��N  �U�U��< t<	t<
t<uB��0�B���/  �$�5�Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �"  =�����.  � 
��`�E�;���  }�ع��E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��K
3��E��EԉE؉E܋E΋��  3�#�#ʁ� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uB�E����u9u�u9u�u3�f�E���  f;�u!B�C���u9su93u�ủuȉu���  �u��}��E�   �E��M���M���~R�DĉE��C�E��E��M��	� �e� ���O��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?�����  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋M��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9M�w�Mԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�B�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�U�f�EċE؉EƋE܉E�f�U��3�f�����e� H%   � ���e� �Ẽ}� �<����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[誘���Ð�.;/�/�/	0A0U0�0�011�0��U���t�p�3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�f��t�C-��C �u�}�f��u/��u+��u'3�f;�����$ f��C�C�C0�S3�@�  ��  f;���   3�@f��   �;�u��t��   @uhL��Qf��t��   �u��u;hD��;�u0��u,h<��CjP蓚����3���tVVVVV�ר�����C�*h4��CjP�g�����3���tVVVVV諨�����C3��q  �ʋ�i�M  �������Ck�M��������3���f�M� 
�ۃ�`�E�f�U�u�}�M�����  }���ۃ�`�E�����  �E�T�˃������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE��P
3ɉM��M��M�M��M��3�� �  �u���  #�#֍4
����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��{����M�����?  ��  f;���  �E�3҉U��U��U�U��U��ɋ�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��V���3�3�f9u���H%   � ���E��\���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �^�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[蒏���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95�*��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��ź��Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��3�PPjPjh   @hT��Dq��	á�	V�5 p���t���tP�֡�	���t���tP��^���������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U���SVW3�jSS�u�]��]������E�#��U���tYjSS�u������#ʃ����tA�u�}+����   ;���   �   Sj�LqP�`p�E���u�w����    �l���� _^[��h �  �u�  YY�E���|
;�r�����P�u��u�:�������t6�+��xӅ�wϋu��u��u��   YY�u�j �LqP�Pp3��   �����8u������    ����u��;�q|;�skS�u�u�u����#�����D����u����YP�Hq�����H��E�#U���u)�����    �������Lp��u�#u��������S�u��u��u�9���#���������3��������U��S�]V�u������@������0�A$�W�y����   ���� @  tP�� �  tB��   t&��   t��   u=�I��
�L1$��⁀���'�I��
�L1$��₀���a��I��
�L1$�!���_^[u� �  ]����% �   @  ]Ë�U��EV3�;�u�s���VVVVV�    �z�����jX�
��3�^]Ë�U����  �ȃ�f9M��   S�u�M������M�Q3�;�u�E�H�f��w�� ���aV�   ��f9u^s)�E�Pj�u����������Et9�M싉�   f����q�M�jQj�MQPR�E�P�*  �� ���Et�E�8]�t�M�ap�[�Ë�U����u�M��h����}�}3���u�u�u�u�q�}� t�M��ap��Ë�U����p�3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[�����Ë�U����u�M��\����E��~�M��Jf�9 t	AA��u���+�H�u �uP�u�u�u�pp�}� t�M��ap����%0p�����̋M�����M�����	���T$�B�J�3��h����H������M�����M����	���T$�B�J�3��:����|��׀���M���q���M������M������M���q���M���q���M������M��|����M��t���j j h8�E�P������ËT$�B�J�3��Ƀ������f����M��q����l����q���M��xq���M������M������M��`q���M������M��Pq����l����Eq����4����:q����P����/q���M��'q���M�������M�������M������M������M������M���p���M������M������M������M������M������M��w����T$�B��0���3��߂�����|���M�������M��I����M��p���T$�B�J�3�謂���(��I���M�����j j h8�EP茖�����j j h8��H���P�s�����ÍM�������M�������E����   �e���M������ÍM������M������T$�B��D���3������L��~���������̍M������M��p����T$�B�J�3������ȱ�~���M������M��E����E����   �e���M�=���ËT$�B�J�3�见�����D~���M��I����M������T$�B�J�3��|����8��~���M������E����   �e���M������ËT$�B�J�3��@����l���}���M�������M������T$�B�J�3���������}���M������M��o����E����   �e���M�n��ËT$�B�J�3��р���ܲ�n}���M�C����T$�B�J�3�讀�����K}���M�� ����T$�B�J�3�苀���4��(}���E����   �e���M�����ÍM�������M�������M��������p���������M��������P��������M������M������M�������`���������@��������M������T$�B��@���3������X��|���M���B���M�����B���M���0��B���M���H�B���M���`�B���M���x�B���M����   �B���M����   �B���T$�B�J�3��r�����|���M��dB���M����YB���M���0�NB���M���H�CB���M���`�8B���M���x�-B���M����   �B���M����   �B���T$�B�J�3���~���H��{���M��n�����|����c���������X�����<����M����M��E����M��=����M��5�����\����*����M��"����M�������L���������l���������,���������������������������������������������������������������M������M�������l���������L��������M������T$�B������3���}������z���������k���������`����������U�����(����J����M��B����������7�����x����,����������!���������������(������������� ����������������x���������H����߿����H����Կ����h����ɿ����X���龿����x���鳿��������騿���M�頿��������长����X���銿����h��������������t����������i����������^����������S���������H����������=����������2����������'�����h��������M������M����������������x�����������������������������������վ���������ʾ�������鿾����8���鴾����X���驾����h���鞾���M�閾���M�鎾����(���郾����H����x�����8����m����������b����������W����������L����������A����������6���������+�����8���� �����X��������M������M����������������������������8��������T$�B��T���3��L{�������w���M�龽����\����i����0�����h���M�頽���M�阽���M�鐽����0�����h���M��}����M��u����M��m����M��e����M��]����M��U����M��M����M��E����M��=����M��5����M��-����M��%�����L���������x��������M������M�������� ���������� �������������޼���M��ּ����<����˼���M��ü����h���鸼���M�鰼���M�騼���M�頼���� ���镼����<���銼����h��������T$�B������3���y���ܷ�v���M�Y�����`����N����M��F����M��>����M��6�����p����+����M��#����M�������P���������4�������������������������������������������ٻ����(����g����D����g���M��g���M��g���M�髻���M�飻���M�電���M�铻���M�鋻���M�郻���M��{����T$�B������3���x��� ��u���M��f���M��M����M��E�����D����f����D����f���M��'����M������M��.���M�������p��������M��������P���������4��������M��޺����`����Ӻ���M��˺���M��ú���T$�B��0���3��+x������t����������e���M�钺���M�銺����(�����e����(�����e����`����i����������e���M��V����M��N�����(����e����(����e���������}e���M��%����M�������(����be����(����We���M�������M�������M������M��'-���M��O-���M��׹���M��Ϲ���M��ǹ���M�鿹���M�鷹���M�鯹���M�駹���M�韹���M�闹�������錹����`���遹��������v����M���,����D����c����M��[����M��S����M��K���������@�����`����5���������*����M��"����M����������������`�������������������������������������������x���������͸���������¸���M�麸���M�鲸���������w�����`���霸���M�锸��������鉸���������~����M��v����M��n����������c����������X���������M����T$�B��D���3��u������Rr����������������̍M������E����   �e���M� ���ËT$�B�J�3��ju�����r�����̋E����   �e���M����ËT$�B�J�3��2u������q�������������̍M阷���M��`����T$�B�J�3���t���L��q���M��=����M��b���T$�B�J�3���t������mq���M��B����M��j����M��"����M��Z����M��R����M��
����M�������M��Zb���T$�B�J�3��ut������q���M������M������M�������M�������M�������M������M������M���a���T$�B�J�3��t�����p���M�錶���M������M��l����M������M������M��T����M��,����M������M��<����M��a���T$�B�J�3��s���l��Lp���M��!����M��I����M������M��9����M��1����M�������M�������M������M�������M��)a���T$�B�J�3��Ds������o����4���鳵����4���騵�������靵�������钵�������釵����$����|�����@����q����� ����f�����0����[��������������T$�B�����3��r���J�3��r���T��Ko���M�� ����T$�B�J�3��r���п�(o���M���9���M���$�B`���M���@�7`���M���\�,`���M����   ������T$�B�J�3��9r�������n���M��9���M��$��_���M��@��_���M��\��_���M���   �����M���   �^����T$�B�J�3���q���@��vn����0����X����������=����������2����������'�������������� ������������������T$�B������3��nq���J�3��dq������n��������������������ȳ����p���齳����`���鲳����(���駳���� ���霳�������鑳����`���醳����p����{���������p����� ����e�����(����Z�����p����O����������D����������9�����D����>�����4����#�����`���������p������������������ ����������(���������`���������p����ֲ��������˲���� ����������(���鵲����p���骲����`���韲����8���锲��������鉲���������~�����8����s����������h����������]����T$�B������3���o���J�3��o������Xl���E���   �e���M����ÍM������M��ܬ���T$�B�J�3��wo���D��l���������f����������[����������������d����ű����T���麱��������鯱����(���餱����D���陱����d���鎱����T���郱���������x�����(����m�����D����b�����l����W����������L�����t����\����t����\���������+�����t���������l����ū���������*�����D����������P����ī����l���陫���������������x����S����T$�B��L���3��;n���J�3��1n���h���j��������頰��������镰��������銰��������������������[���������[���������^����������S����������[���������[���������B����������'����������������������������������������������d������������������������گ����d����ϯ���������į��������鹯��������鮯����t���飯��������阯����T���鍯����D���邯���T$�B������3���l���J�3���l���l��}i�����������̋M��H����M���L�=����M���\�2����M���p�'����T$�B�J�3��l������/i�������������̋M�������M���L�����M���\�����M���p�׮���T$�B�J�3��Bl�������h�������������̋M����c���T$�B�J�3��l���L��h�����������̋M���H�%����T$�B�J�3���k���x��}h�����������̋T$�B�J�3��k������Xh������̋EP�M�Q������ËT$�B�J�3��k���d��'h�����̋M������T$�B�J�3��ck������ h��������������̋EP�M�Q胿����ËT$�B�J�3��*k�������g�����̋M��^���M����]����M��� �R����M���<�G����M���X�<����T$�B�J�3���j�����tg��̋M��R^���M��������M��� �����M���<������M���X�����T$�B�J�3��j���`��$g��̍M��ȧ���T$�B�J�3��cj���J�3��Yj�������f����̍M�阧���T$�B�J�3��3j���J�3��)j�������f����̋M��Ty���T$�B�J�3��j�����f��������������̋EP��|��YËE����   �e���M�����ËT$�B��\���3��i���H��Qf���������������̍M������T$�B�J�3��i���J�3��yi���t��f����̍M�鸦���T$�B�J�3��Si�������e��������������̋E�P�7|��YËE����   �e���M��m���ËT$�B��\���3��i���l��e���������������̋EP�M�Q�#�����ËT$�B�J�3���h������ge�����̍M������M�� �����l���������T$�B��t���3��h�����*e��������̋M��w���T$�B�J�3��ch������ e��������������̋M��ؐ���T$�B�J�3��3h�������d��������������̍M���-���T$�B�J�3��h������d��������������̋T$�B��l���3���g���J�3���g���H��kd���������̍�L����ņ��������麆���T$�B������3��g������/d�������������̍M��[���T$�B�J�3��cg���8�� d��������������̋EP�M�Q胻����ËT$�B�J�3��*g�������c�����̋M��؝���T$�B�J�3��g������c��������������̋M���P�����T$�B�J�3���f������mc�����������̍M�ȅ���T$�B�J�3��f�����@c��������������̍M�X,���T$�B�J�3��sf���H��c��������������̍M�騣���E�P�M�Q苺����ËT$�B�J�3��2f���J�3��(f�������b���̍M��+���T$�B�J�3��f������b��������������̋M��X����T$�B�J�3���e���T��pb��������������̋E����   �e���M��X�ł��ËM���ɂ���T$�B�J�3��e������!b���������������̋E����   �e���M��P�u���ËM���y����T$�B�J�3��4e�������a���������������̍M�鈍���T$�B�J�3��e�����a��������������̍M��X����M��*���T$�B�J�3���d������ha������̍M������M�� ����T$�B�J�3��d���J�3��d�����.a������������̋M����š���T$�B�J�3��`d�������`�����������̍M,�����M�����T$�B�J�3��+d�������`������̍M,鸥���M鰥���M�騥���T$�B�J�3���c������`��������������̋M�������T$�B�J�3���c���(��``���������������j j h8�E�P�w����ËM������T$�B�J�3��}c���\��`���M���V���T$�B�J�3��Zc�������_���M��)���T$�B�J�3��7c�������_���M���(���M����n����T$�B�J�3��	c������_���M��V���u���u��YËT$�B�J�3���b�����y_���M������T$�B�J�3��b���X��V_���T$�B�J�3��b���@��;_����������h�k����Yù��U��h�k����Y�h�k�����YùX�`U��h�k����Y�h�k�ڇ��YÃ= uK���t���Q<P�B�Ѓ��    ���tV����O��V��N�����    ^ù��U�����'���X�U���Y�#]��   �� �� �� �� �� � 4� L� T� p� �� �� �� �� �� �� � &� :� L� \� h� v� �� �� �� �� �� �� �� � � (� 6� B� P� Z� j� t� �� �� �� �� �� �� �� ��  � � � 0� <� L� ^� r� ~� �� �� �� �� ��  � � 4� D� Z� t� �� �� �� �� �� �� �� � *� @� P� `� p� �� �� �� ��     ��         <k^ktk0kRk        ���2t5�CV        �B�V                    %LM       �   �� �� bad allocation  <��! � ` ��0 ��� P �a3D-COAT Start import!   To import a new object? File exists!    export.txt  Folder ..\MyDocuments\3D-CoatV3\Exchange not found! 3D-CoatV3   Exchange    preference.ini  3D-Coat.exe is run! 3D-Coat.exe not found!  open    
             �?]   autopo  curv    prim    alpha   vox retopo  ref uv  ptex    mv  ppp [   # end   v       # begin      vertices
            �?vt   texture vertices
  /   f   usemtl   faces
 g   mtllib  mtl map_    illum 2
    Tr 0.000000
    Ns 50.000000
   Ks  Kd  Ka 0.300000 0.300000 0.300000
  newmtl  No selected objects!    Object "    " has no UVW tag.
UV coordinates can't be exported. Material not found on   object. Default Name    Export object   #Cinema4D Version:  %d.%m.%Y  %H:%M:%S  #File created:  #Wavefront OBJ Export for 3D-Coat
  File     write success!   ��import.txt  output.obj  obj ��`� �<��� ��p� ��p� t�p� ���� `� @� �� �� �� ��  � p� `� ��           Y@إ�� �� �� �� �� � �� �@� `� �� �� ��  � � ��� �� �� � �� �@� �� �� �� �� l��� �  �  � �� �� �� �� Selection   Error on inserting phongTag. Object:    Create objects...   Memory allocation error for material.   ��@� -���� 0��� �"�"���7`�����������H���vector<T> too long  bad cast    ios_base::eofbit set    ios_base::failbit set   ios_base::badbit set    �� =    X       P   f   vt  Gathering of data...     not found!  can not removed!   normalmap   displacement %f displacement    map_Ks %s   map_Ks  map_Kd %s   map_Kd  Ke %lf %lf %lf  Ke  Ks %lf %lf %lf  Ks  Ka %lf %lf %lf  Ka  Kd %lf %lf %lf  Kd  illum %d    illum   d %lf   d   Ns %lf  Ns  newmtl %s    open!  vt %lf %lf %lf  vt %lf %lf  v %lf %lf %lf   g %s    mtllib %s   Parse file...   Open file:  .   textures.txt    \��Q�OP� �`��0� �icon_coat.tif        �f@-DT�!	@���`�p������������a     @�@���`�p��������������@� �0���К@����������T��`�p����������������`�p������������� �0�@�P�`�p�����Ц�����~   %s      B   KB  MB       P? GB     ����MbP?$� a0Gl��`�� e �0�cК@�0c������d          �#   M_EDITOR    ���res    ? �Ngm��C   O�������^            ���*   C   ����d����string too long invalid string position r            
   !   "   2   *            #   3   +       w   a   r b     w b     a b     r +     w +     a +     r + b   w + b   a + b   ����;�����                  �?      �?3      3            �      0C       �       ��                    �?      �?3      3                      �                     ���e��Unknown exception   ����csm�               �                                                                                                                                                                                                                                                                                                      ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������LC_TIME LC_NUMERIC  LC_MONETARY LC_CTYPE    LC_COLLATE  LC_ALL  p�    o�d���o�X�����L�����@���Q�8�����	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ _., _   ;   =   =;  |\���bad exception   EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    ��e+000          �~PA   ���GAIsProcessorFeaturePresent   KERNEL32          �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:    ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx                      �������             ��      �@      �              �?5�h!���>@�������             ��      �@      �        HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun united-states   united-kingdom  trinidad & tobago   south-korea south-africa    south korea south africa    slovak  puerto-rico pr-china    pr china    nz  new-zealand hong-kong   holland great britain   england czech   china   britain america usa us  uk  swiss   swedish-finland spanish-venezuela   spanish-uruguay spanish-puerto rico spanish-peru    spanish-paraguay    spanish-panama  spanish-nicaragua   spanish-modern  spanish-mexican spanish-honduras    spanish-guatemala   spanish-el salvador spanish-ecuador spanish-dominican republic  spanish-costa rica  spanish-colombia    spanish-chile   spanish-bolivia spanish-argentina   portuguese-brazilian    norwegian-nynorsk   norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg   german-lichtenstein german-austrian french-swiss    french-luxembourg   french-canadian french-belgian  english-usa english-us  english-uk  english-trinidad y tobago   english-south africa    english-nz  english-jamaica english-ire english-caribbean   english-can english-belize  english-aus english-american    dutch-belgian   chinese-traditional chinese-singapore   chinese-simplified  chinese-hongkong    chinese chi chh canadian    belgian australian  american-english    american english    american    l�ENU X�ENU D�ENU 8�ENA 0�NLB $�ENC  �ZHH �ZHI �CHS  �ZHH �CHS ؔZHI ĔCHT ��NLB ��ENU ��ENA ��ENL x�ENC d�ENB X�ENI H�ENJ <�ENZ $�ENS �ENT ��ENG �ENU �ENU ԓFRB ēFRC ��FRL ��FRS ��DEA |�DEC h�DEL X�DES H�ENI 8�ITS ,�NOR �NOR �NON �PTB ؒESS ȒESB ��ESL ��ESO ��ESC t�ESD d�ESF P�ESE <�ESG (�ESH �ESM �ESN ��ESI �ESA БESZ ��ESR ��ESU ��ESY ��ESV x�SVF p�DES l�ENG h�ENU d�ENU \�USA T�GBR L�CHN D�CZE <�GBR ,�GBR $�NLD �HKG �NZL �NZL ��CHN �CHN �PRI ܐSVK ̐ZAF ��KOR ��ZAF ��KOR ��TTO l�GBR ��GBR p�USA h�USA 6-0   OCP ACP Norwegian-Nynorsk   c c s   U T F - 8   U T F - 1 6 L E     U N I C O D E    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   %   ->* &   +   -   --  ++  ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(    $���������؝̝���r�������������L�����������������P{����|�x�t�p��sl�h�d�`�\�X�T��zP�L�H�D�@�<�8�4�0�,�(�$� �������؜̜����x�X�8����؛����l�P�@�<�4�$� ����ܚ����x�P�(���������l�@�$��r_nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp       SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    1#QNAN  1#INF   1#IND   1#SNAN  CONOUT$     H                                                           p���^   RSDSF]I(.�L���,8�eU   C:\Program Files\MAXON\CINEMA4D_Architecture_Edition_R11010\plugins\AppLink_3DCoat\obj\Applink_3DCoatR11_Win32_Release.pdb              �P�           `�l���    �       ����    @   P� �        ����    @   ��           ����                @�Т           ���    @�       ����    @   Т\�        ����    @   $�           4��                x�P�           `�h�    x�        ����    @   P�           ����h�    ��       ����    @   ��           ̣أh�    ��       ����    @   ��            ���           �$�@�    ��       ����    @   ���       ����    @   \�           l�t�    ��        ����    @   \�           ���           ��Ȥ�<�X�    �       ����    @   ��L�              P    �           � �$�@�    L�       ����    @    ���              @   ���              @   \�            L� �            ����           ����أh�    ��       ����    @   ��            ���           ���    ��        ����    @   �            ��4�           D�P��    ��       ����    @   4�            0���           ������h�    0�       ����    @   ��    P       P�Ц           ���Ȥ�<�X�    P�       ����    @   Ц            ��(�           8�D��    ��       ����    @   (�            ��t�           �����    ��       ����    @   t�             ���           Чܧ�     �       ����    @   ��             ��           �,����     �       ����    @   �            @�\�           l�|�ܧ�    @�       ����    @   \�    X       ����           ��ԨȤ�<�X�    ��       ����    @   ��            ��(�    ��       ����    @   ���        ����    @   D�           T�(�                ��p�           �����(�    ��       ����    @   p�             ���            (�ԩ           ����    (�       ����    @   ԩ            D� �           0�8�    D�        ����    @    �            `�h�           x�����    `�       ����    @   h�            x���           ĪԪ����    x�       ����    @   ��            ��    ��        ����    @   �            ��8�           H�P�    ��        ����    @   8�            ����           �����    ��       ����    @   ��            �̫           ܫ�8�    �       ����    @   ̫            ��D�            t�,�           <�H�h�    t�       ����    @   ,�            ��x�           �������    ��       ����    @   x�            |�Ȭ           ج�    |�        ����    @   Ȭ            \�$�            d�$�           4�@��    d�       ����    @   $�            4�p�           �����    4�       ����    @   p�        �� �� pT �� � CI qI �I �J �J �K �K L /L kL �L �L �L  M �M 9N �N �O \R �S �T }U �W AX yX �X �X 6Y �Y �Y gZ �Z  [ r[ �[ :\ �] 4^ m_ �` a ia �a �a �a !b Hb �b �b $c Hc xc �c �c (d Xd �d �d e He xe �e �e f Hf �f �f �f g 8g yg �g �g 'h wh �h �h i Ki �i �i �i .j Qj tj �j �j �j k                 ����0I    8I"�   8�                       ����^I    fI"�   l�                       "�	   į                       �����I    �I   �I   �I    �I    �I    �I    �I    �I"�   0�                       �����I    J   J����J    J   (J   0J   8J   @J   KJ	   VJ
   aJ	   aJ   aJ   aJ   aJ   iJ   qJ   yJ   �J   �J   �J   �J   �J   �J   �J   �J   �J�����J    �J   �J"�   �                       "�	   p�                       ����8K����QK   YK����YK   aK   zK   �K����K����"K�����K    �K"�   ��                       �����K    �K   �K"�   �                       ����L    'L"�   (�                       ����JL    RL"�   \�                       �����L    �L"�   ��                       �����L    �L   �L"�   Ĳ                       �����L"�    �                       ����M"�   ,�                       "�   |�                       ����;M    TM    \M    dM    lM    wM    M    �M    �M    �M    �M    �M    �M"�   �                       �����M    �M   �M   �M   N   N   N   +N"�   l�                       ����TN    \N   gN   rN   }N   �N   �N   �N"�   д                       �����N    �N   �N   �N   �N   �N   �N    �N�����N   �N	   O
   O   O   O   &O   1O   <O   GO   RO   ]O   hO   sO   ~O   �O   �O   �O   �O"�B   ̵                       �����O    �O   �O   �O   �O   �O   �O    �O�����O   �O	   	P
   P   P   *P   5P   @P   KP   VP   aP   lP   wP   �P   �P   �P   �P   �P   �P   �P   �P   �P   �P   �P   �P    Q!   Q   Q#   $Q$   ,Q%   4Q&   ?Q'   JQ(   UQ)   `Q*   kQ+   vQ,   �Q-   �Q.   �Q   �Q0   �Q1   �Q2   �Q3   �Q4   �Q5   �Q6   �Q7   �Q8   �Q9   
R:   R;    R   +R=   3R>   ;R?   FR@   QR"�$    �                       ����zR    �R   �R   �R   �R   �R   �R   �R   �R   �R    �R
   �R   �R   �R    �R   �R   S   S   S    S   &S   1S   9S   AS   LS   WS   bS   jS   uS   }S   �S   �S   �S    �S!   �S"   �S"�   D�                       �����S    �S   �S    �S   �S   T   
T   T   T   %T	   0T
   ;T   FT   QT   \T   gT   rT   }T   �T   �T   �T   �T   �T   �T   �T   �T"�   8�                       �����T    �T   �T   �T    U    U    U    !U   )U   1U	   <U
   DU   OU   ZU   bU   mU   uU"�?   �                       �����U    �U   �U   �U    �U    �U    �U   �U   �U   �U   �U   V   V   V   #V   .V   9V   AV   IV   QV   YV   aV   iV   qV   yV   �V   �V   �V   �V   �V   �V   �V   �V   �V!   �V"   �V"   �V$   �V%   �V&    W'   W"   W)   W*   &W+   1W,   <W"   GW.   RW"   ]W0   hW1   sW0   �W3   �W4   �W5   �W0   ~W0   �W0   �W0   �W:   �W;   �W<   �W   �W����(X     X"�   ܼ                       ����`X"�   �                       �����X    �X"�   <�                       �����X    �X"�   p�                       "�   Ƚ                       �����X�����X   Y   Y   Y   Y   &Y   .Y"�   ,�                       ����QY����YY   aY   iY   qY   yY   �Y   �Y"�
   ��                       �����Y�����Y   �Y   �Y   �Y   �Y   �Y   �Y   �Y   �Y"�
   �                       ����Z����Z   'Z   /Z   7Z   ?Z   GZ   OZ   WZ   _Z"�
   x�                       �����Z�����Z�����Z�����Z   �Z�����Z   �Z   �Z   �Z�����Z����["�   ȿ                       "�   �                       ����;[    C[   N[   Y[   d["�   d�                       �����[    �[   �[   �[   �[   �["�   ��                       �����[    �[   \   \   \   $\    /\"�#   �                       ����b\    m\   x\   �\   �\   �\   �\   �\   �\   �\	   �\
   �\   �\   �\   �\   ]   ]   ]   (]   3]   >]   I]   T]   _]   j]   u]   �]   �]   �]   �]   �]   �]   �]    �]!   �]����^    $^    ,^"�   ,�                       "�   ��                       ����O^    Z^   e^   p^   {^   �^   �^   �^   �^   �^	   �^
   �^   �^   �^   �^   �^   �^   
_   _    _    _   +_   6_   A_   L_   L_   W_   b_"�   ��                       �����_    �_�����_   �_   �_�����_�����_   �_   �_�����_����`
   `
   `   $`   /`   :`   E`
   P`   [`   f`   q`   |`
   �`   �`   �`   �`   �`�����`    �`   a   a"�   h�                       ����@a    Ha   Sa   ^a"�   ��                           P�      �   �(�    @�    ����       `�     \�    ����       �������a"�   D�                       �����a"�   p�                       @           �@           	����    ����                  "�   ��    �                           ��              ��@           �
             (�����        b����    "�   L�   8�               ����@b"�   ��                       @           \             ������        pb����    "�   ��   ��               "�   8�                       �����b    �b   �b   �b   �b"�   ��                       �����b    �b   c   c   c����@c"�   ��                       ����pc"�   ��                       �����c"�   �                       �����c    �c�����c"�   0�                       ���� d"�   l�                           p    ��   ����(�     �    ����    (    &    ��    ����    (    %����Pd"�   ��                           Z�    ,�   8�(�    d�    ����       =������d    �d�����d"�   T�                       @           �)             ������        �d����    "�   ��   ��                   @    <����� e����e����e"�    �                          L�h�(�    @�    ����    (   �+     �    ����    (   +����@e"�   ��                       ����pe"�   ��                       �����e"�   ��                       @           �/@           �/����    ����    ����    ����    "�   (�   l�                             �            �@           �3@           �2"�    �   ��                             ��            ������    ����    ���� f              ����f����@f"�   0�                       @           �6             \�����        pf����    "�   ��   l�               �����f"�   ��                       �����f"�   ��                       ���� g"�   �                       ����0g"�   @�                       @           �;            l�����`g           hg        "�   ��   |�               @           �>            ��"�   �   ��               �����g����    ����                         �����g"�   L�                       ���� h            h"�   x�                       ����Ph            lh"�   ��                       @           >D            ��"�   8�    �               �����h                                     @           	F            h�"�   ��   x�               �����h    �h                                     @           �J@           �I"�   T�   ,�                             ��            ������    ����    ���� i              ����i����@i"�   ��                       ����pi    xi"�   ��                       �����i    �i   �i"�   ��                       �����i"�    �                       ����j����&j"�   L�                       ����Ij"�   ��                       ����lj"�   ��                       �����j    �j"�   ��                       �����j    �j"�   �                           ��    |������j"�   P�                          ����(�    ��    ����    (   ������    ����    ����    I�    ����    ����    ����    z�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    u�        A�����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    /�    ����    ����    ����    f�    ����    ����    ������    ����    ����    ����    ��    ����    ����    ����    R�    ����    ����    ����    ~    ����    ����    ����    �        �        �    ����    ����    ����    �    ����    ����    ����        ������    ����    ������@           �����    ����                  �"�   �   ,�                   ����    ����    ����    �    NW����    ����    ������    ����    ����    ����^b    |    ��   ��(�    4�    ����       "    ����    ����    ����    M%����    \%����    ����    ����    '����    '����    ����    ����B)F)    ����    ����    �����)�)    ����    ����    ����    y+    ����    ����    ����    �.    ����    ����    ����    �2    ����    ����    �����4�4    ����    ����    ����    I    ����    ����    ����[[    ����    ����    ����    be    ����    ����    ����    Cf    ����    ����    ����    
j    ����    ����    ����    [k    ����    ����    ����    �m    ����    ����    ����    Lo    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    y�    ����    ����    ����    ��    ����    ����    ����    @�    ����    ����    ��������    ����    ����    ����Q�h�    ����    ����    ��������    ����    ����    ����    s�    ����    ����    ����    1    ����    ����    ����    �    ����    ����    ����    C    ����    ����    ����    	        E����    ����    ����    !!8�         ��  p ��         � Tq                     �� �� �� �� �� � 4� L� T� p� �� �� �� �� �� �� � &� :� L� \� h� v� �� �� �� �� �� �� �� � � (� 6� B� P� Z� j� t� �� �� �� �� �� �� �� ��  � � � 0� <� L� ^� r� ~� �� �� �� �� ��  � � 4� D� Z� t� �� �� �� �� �� �� �� � *� @� P� `� p� �� �� �� ��     ��     C CloseHandle EProcess32Next Module32First CProcess32First  � CreateToolhelp32Snapshot  KERNEL32.dll  ShellExecuteExA SHELL32.dll �InterlockedIncrement  �InterlockedDecrement  !Sleep �InitializeCriticalSection � DeleteCriticalSection � EnterCriticalSection  �LeaveCriticalSection  �RtlUnwind -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent ZRaiseException  �GetLastError  �HeapFree  � DeleteFileA �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �LCMapStringA  zWideCharToMultiByte MultiByteToWideChar �LCMapStringW  [GetCPInfo �GetModuleHandleW   GetProcAddress  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �SetLastError  RGetACP  GetOEMCP  �IsValidCodePage �GetModuleHandleA  �HeapCreate  �HeapDestroy WVirtualFree TVirtualAlloc  �HeapReAlloc �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA �WriteFile �GetConsoleCP  �GetConsoleMode  AFlushFileBuffers  hReadFile  �SetFilePointer  ExitProcess �GetModuleFileNameA  JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW �GetEnvironmentStringsW  TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �HeapSize  �GetLocaleInfoA  =GetStringTypeA  @GetStringTypeW  mGetUserDefaultLCID  � EnumSystemLocalesA  �IsValidLocale �InitializeCriticalSectionAndSpinCount �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW �SetStdHandle  �LoadLibraryA  �GetLocaleInfoW   CreateFileW x CreateFileA �SetEndOfFile  #GetProcessHeap      %LM    ��          �� �� �� �� �   Applink_3DCoatR11.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �q$|    .?AVApplinkDialog@@ $|    .?AVGeDialog@@  �q�q$|    .?AVbad_alloc@std@@ $|    .?AVexception@std@@ $|    .?AVfacet@locale@std@@  $|    .?AVcodecvt_base@std@@  $|    .?AUctype_base@std@@    $|    .?AVios_base@std@@  $|    .?AV?$_Iosb@H@std@@ $|    .?AV?$basic_istream@DU?$char_traits@D@std@@@std@@   $|    .?AV?$basic_ios@DU?$char_traits@D@std@@@std@@   $|    .?AV?$ctype@D@std@@ $|    .?AV?$basic_streambuf@DU?$char_traits@D@std@@@std@@     $|    .?AV?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    $|    .?AV?$codecvt@DDH@std@@ $|    .?AV?$basic_istringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    $|    .?AV?$basic_filebuf@DU?$char_traits@D@std@@@std@@   $|    .?AVlogic_error@std@@   $|    .?AVruntime_error@std@@ $|    .?AVlength_error@std@@  $|    .?AVfailure@ios_base@std@@  $|    .?AVbad_cast@std@@  $|    .?AV?$basic_ifstream@DU?$char_traits@D@std@@@std@@  �q�q$|    .?AVCommandData@@   $|    .?AVBaseData@@  $|    .?AVApplinkPreferences@@    �q�q�q$|    .?AVGeModalDialog@@ $|    .?AVGeUserArea@@    $|    .?AVSubDialog@@ $|    .?AViCustomGui@@    �q�q�q�q�q�q�q�q�q$|    .?AVGeSortAndSearch@@   $|    .?AVNeighbor@@  $|    .?AVDisjointNgonMesh@@  �q$|    .?AVTexturePreview@@    �q�q�q�q�q�q�q�q�q�q�q�q�q�q�����q$|    .?AV_Locimp@locale@std@@    �q   �q$|    .?AVout_of_range@std@@  �q�{�{�{�{�{�{�{�{�{�{ ||||        �q
   Copyright (c) 1992-2004 by P.J. Plauger, licensed by Dinkumware, Ltd. ALL RIGHTS RESERVED.      N�@���D�q$|    .?AVtype_info@@             u�  s�          �q            fmod         ��Ơ_�Ơ$�Ơ_�Ơ]�]���]�ƠƠ_�Ơsqrt    0~2�   4�        �q$|    .?AVbad_exception@std@@ ��������    �q                                                                                                                                                                                                                                                                                                                                                abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     p��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����    C                                                                                              ��            ��            ��            ��            ��                              @        0~��8����   ��p�                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                         ?�?�?�?�?�?�?�?�?�?�?  ?                                                                                                                                                                                                                                                                                           `    `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����
                                                          ׄ      x   
          ��   ��	   `�
   Ȍ   ��   l�   H�   �   �   ��   ��   L�   $�   �   ��    h�!   p�"   Јx   ��y   ��z   ���   ���   ��\�L�       ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      ������%�*�0�6�<�B�^�c�y�~�������΢����2�F�^�r���������֣���6�;�U�Z�z�������ڤߤ�����2�J�^�~�������¥֥��"�'�A�F�f�z���  l�h�d�`�\�X�T�L�D�<�0�$������ �������������؏̏ď����������������x�t�p�d�P�D�	         �.   <���������@   .       �            �&         ��   �   ԇ   ؇    �   �!   �   ̇   ć   ��   �    �   ��   ��    ��   ��   ��   ��   ��   �   �   ��   ؟   П"   ̟#   ȟ$   ğ%   ��&   ��      �      ���������              �       �D        � 0                                                                                                                                                                                                                        �p     ����    PST                                                             PDT                                                             � 	����        ����           ���5      @   �  �   ����             ������������   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l           �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                                                                                                                                                                                       �   00A0V0d0�0�0�0�0:1$2M2�2�2�2@3V3m3�3�3�3�344&4>4b4}4�4f6{6�6h7�7�7�7�7�8�8�89l9�9	:c:�:�:�:;0;}<�<�<V=g=�=6>K>�>�>�>�>�>f?�?�?�?      �   	0A0m00�0�011'1>1Y1q12D2U2q2�4�4�45&5>5r5�5�5,6A6U6e6�6�6�6�6�6�6R7g7�7�7�7?8l8�8�8�89^9�9�9�9Z:}:�:�:�:; ;7;;�;�;�;�;�;<<4<u<=*=@=T=b=�=�=�=�=�=>'>M>j>�>�>�>�>?7?W?n?�?�?�?�? 0  �    000/0B0p0t0x0|0�0�0�0�0�0�0�0�0�0�2�2F4[4q4�4�4�4�4�4515I5b5{5�5�5�5�5�5
66%6>6S6[6q6�6�7�7�7�7�78838L8e8}8�8�8�8�8�8+9=9O9X9m99�9�9�9:#:9:O:j:�:�:�:�:;;$;?;T;�;�;�;�;	<$<N<c<x<�<�<�<�<�<�<�<==B>X>q>�>�>�>�>�>??9?R?k?�?�?�?�?�?   @    00%010?0X0m0v0�0�0�1�1�12%2>2W2o2�2�2�2�2�23)3:3W3l3�3�3�3�3�3�3�3�344:5P5i5�5�5�5�5�5�5616J6`6u6�6�6�6�6�677.767O7d7m7�7�7�8�8�89959N9f99�9�9�9�9�9:.:e:v:�:�:�:�:;;2;O;c;y;�;�;�;<<.<l<�<�<=!=7=I=[=c=y=�=�=�=>">I>_>�>�>�>�>�>�>??+?c?y?�?�?�?�?�?   P  $  70H0Z0c0y0�0�0�0�01#191O1l1�1�1�1�1�1�1=2U2j2�2�2�2�2�2�2#393R3k3�3�3�3�3�344$4@4�4�4�4�4�4�45&5=5o5�5�5�5�5�5�56+6e6w6�6�6�6�6�6�6+7=7O7X7m77�7�7�78)8?8U8p8�8�8�899.9J9_9�9�9�9�9�9�9::$:9:;*;>;V;o;�;�;�;�;�;�;<.<G<b<==0=9=N=`=�=�=�=�=�=�=>#>U>k>>�>�>�>�>?,?f?{?�?�? `  �   0V0h0z0�0�0_1s1�1�1�1�1�1�1232L2e2z2�2�2�2�2�2�23,3F3t3�3�3�3�3�34/4D4M4i4�4�4�4�4�4�45555R5d5v5~5�5�5�5�5v6�6�687N7�7�7�7�7
8l8�8�8�8=9S9k9�9�9:A:�:�:(;�;�;�;<P<f<�<�<�<=>=M=�=�=�=�=>�>�>�>�>G?U?s?�?�?�?   p  t   
0 0X0f0w0�0�0�01,1�1�1�1�122#2W2p2�2�2�2�233F3�34R4o45:5U5�5�5�5�5�5�5�6�6�6(7D7c7}7F<�<�>E?�?�?�?�? �  T   0$090d0�0�0,1=1N1W1m1~1�1�1�122>2t2�2�2�2�2	3�394�4�5�78k9�:';2<�=>E?   �  �   T0f0�061F1^1p1�1�1�1�1�1R2h2�3�3y4�4�4�4!5T5�5�56B6d6�6�6�6�668H8^8p8�8�8�89�9�9:�:;;.;@;S;�;�;�;U<r<�<p=�=�=�=�=>F>j>�>?-?�?�?   �  �   0�0�0�0�01"1f1�1�102M2�23�3�3�3!4�4�4�4�4n5�5�5F6f6�6�6�6�6�9.:[:p:�:�:�:�:;!;5;�;�;5<U<�<�<�<%=>=W=p=�=�=>V>�>�>? �  �   60H01j1�1�1�12F2U2�2&383O3f4x4�45"5*5C5X5a5y5�5�56686q6�6�6�6�6*7�7�79�;�;<G<b<{<�<==!=9=N=�=�=�=�=>!>Z>o>�>�>�>�>�>'?@?X?u?�? �  �   	0\0h0}0�0�0D1b1�1�1:2a2}2�2&3V3�3�3x4�4!5?5�5�56�6�6�6?7Z7o7w7�7�7�78.8G8`8x8�8�899#9<9Q9�9�9�9�9:�:�:;%;�;�;)<><�<�<�<#=8=�=�=G>�>???8?L?U?m?�?�?�?   �  �   0+0G0w0�01(162H2�2�23343H3Q3i3�3�3�34'4]4�4�4�4�4�4�4�45c5{5�5�5�5�56 636K6�6�6q7�79919P9�9�:�:�:;S;o;�;<F<l<�<�>�?   �  �   (0�0J1�1f2x2�23383S3�3�3�3,4�4�4�4%5E5�5�5�5�5�56h6�6�6�6�6�6717:7R7f7�7�7�78 8�8�8�8�8	99&9>9�9�9�9�9:�:�:�:<<*<j<x<�<�<�<�<�<=,=A=W=??,?:?�?�?�?�? �  T   00)0B0�1�1�1�1I2T2q2�2�2
3&3<34�56Y6H7h7�89s9�9E:�:�:�:	;;�<�<�=�=�=     8   62E2b2t2�2�2�68(8�8F:X:�:U;�;�;�;�<=�=>>�>�>  0   �2�2f6u6g:�:�:;a;u;�;�;�;f<{<E=�=�>�>     t   �2�35&555\5�5�5�5�5�56&686T6[6w66�6�6�6�6�67�7�7	8F9X9::Q:q:|:�:�:�:�:�:�:;%;L;�;6<D<�<�<�<�<6=H=F>X> 0 P   1+1�4�4�4�4�4�45
55m5z5�566H6�6�6F7T7q7�7�799&:5:�:f;u;^<5=f=x=�>   @ P   F0T01191@1V1�1�1�12292@2V2�2�2�2j4�4�45668E8�;�;�=�=�>�>d?�?�?�?�?   P �   0$090t0�0�0�01*1V1d1�1�1�1�1�12!2D2d2�2�2�2�23$3T3�3�3�34$4Q4a4�4�4�4�45$5I5d5�5�5�5�5$6N6t6�6�6�6�67D7�7�7�748U8f8�8�8�8�8�8�8�8$9^9�9�9�94:T:�:�:�:;4;k;�;�;�;�;<4<T<t<�<�<�<$=D=Z=�=�=�=>D>t>�>�>�>?1?�?   ` t   0�0(1]1�2�2�2�23!3D3q3�3�3�3H4�4�4�4:5\5�5�5�56,6{6�67@7p7�7�8�8�9�9n;�;�;u<}<�<N=�=�=+>g>�>�>?L?�?�?   p T   V0�0�01t3�3�3/4�45�6�6�6*7J798�8�8#9s9�9:s:�:3;�;�;3<�<�<S=�=>s>�>3?�?�? � �   C0�0	1y1�12c2�2�2*3P3�3�3�34>4�4�4�4+535d5�5�56Z6�6�6N7�7�78D8�8�8�8!9T9�9�9:A:q:�:;1;�;�;�;�;<"<�<�=6>�>�>�>�>�>�>�>�>�>�>�?�?�?�?�?�?�? � �    000�0�0�0�0121N1q1�1�1�1�12D2t2�2�2�23T3�3�3�34e44�4$5D5d5�5�5�56D6t6�6�67A7a7�7�78`8�8�8�899d9�9�9:D:^:;4;�;9<�=�=>>%>:>X>b>�>$?D?d?�?�?�?�?�?   � `   s0�0E1�1�1�1$2T2�2�2�2d4�4�45H5M5Y5�5�5{9�9�9�9�9#:M:t:�:�<�<�<�<�<==1=K=_=q=�=�=�=   � �   >146M6v6�6�6�6�6�6:7o7�7�89L9S9�9�9:#:F:d:�:�:�:�:;;4;E;d;u;�;�;�;�;<A<d<y<�<�<�<�<�<=$=D=d=�=�=�=�=>4>T>�>�>�>�>?$?Q?d?�?�?�?   � �   040T0�0�0�0�01$1D1d1�1�1�1�12$2G2}2�2�2�2�23d3�3�3�3�3$4A4t4�4�4�455646T6t6�6�6�6�67A7Q7d7�7�7�7�7�78#818@8a8�8�8�8�8919A9Q9d9�9�9�9�9�9::D:d:�:�:�:�:;$;D;d;�;�;�;�;�;�;$<7<P<_<�<�<�<�<�<1=D=t=�=�=�=>$>D>d>�>�>�>�>?$?D?d?�?�?�?�? � �   0$0T0�0�0�0 1$1D1d1�1�1�1�1242d2�2�2�2�23$3D3d3�3�3�3�3444T4t4�4�4�4515T5t5�5�5�5�56$696P6_6�6�6�6�6�6$7T77�7�78D8h8�8�9�9�9�9�9:_:�:�:�:�:;!;=;h;�;�;�;�;�;<D<�<�<I=e=�=�=I>e>�>�>U?�?�? � �   =0U0�0�01(1L1h1�1�1�1�12(2L2h2�2�2�2�2�2$3D3d3�3�3�3�3�3!4D4t4�4�4�4�4515D5�5�5�5�56!6D6d6�6�6�67$7Q7t7�7�7848T8t8�8�8�8�8949T9q9�9�9�9�9:n:�:�:;G;�;�;!<�<�<�<X=z=�=>.>F>�>�>�>s?�?�?�?   � �   0D0�0�01�1�1�1S2|2�23.3C3�3,4W4�4�415W5�5�516�67<7Y7�7�78~8�8�89a9�9<:d:�:�:�:�:�:;+;P;t;�;�;<1<T<t<�<�<�<=7=�=�=�=>&>:>Y>�>�>�>?$?A?d?�?   �   0#0(0-0I0q0�0�0�0�0111T1�1�1�1242T2q2�2�2�2(3g3�3�34A4T4�4�4�4�4$5D5d5�5�5�5�56616D6a6q6�6�6�6�67A7Q7d7�7�7�78!818A8T8t8�8�8�8�89?9d9�9�9�9�9�9:4:_:�:�:�:�:;D;d;�;�;�;�;<$<D<d<�<�<�<�<=D=�=�=�=C>�>�>�>?D?q?�?�?�?�?  �   0!040T0t0�0�0�0	11r1�1�1�12$2D2�2�2�2�2�2323F3V3�3�3�3�34H4_4w4�4�4�4�45:5X5m5�5�5�5�5�56"626T6�6�6�6;7M7a7q7�7�7848�8�8�8�89/9T9t9�9�9�9�9:$:D:a:t:�:�:�:;4;T;�;�;�;<!<4<d<�<�<�<�<�<�<=�=>2>e>�>�>?e?�?�?�?   �   50u0�01O1�1�12B2u2�23R3�3�34E4u4�4�4%5U5�5�556u6�6�67@7T7d7�7�78U8�8�8%9e9�9�9:9:C:m:r:�:�:�:;);e;�;�;�;E<i<�<�<�<&=O=�=�=�=>V>�>?'?D?d?�?�?�?�?   0 �   00$0A0Q0d0�0�0�0�0�0111Q1t1�1�1�12$2D2d2�2�2�233$3D3d3�3�3�3�344D4o4�4�4�45 5A5T5t5�5�5�5�546G6b6r6�6�6�6�67(7G7�7�7�788A8s8�8�8�8�8�8959G9t9�9�9�9:4:a:�:�:�:;$;D;�;�;�;<4<a<�<�<�<�<=!=D=d=�=�=�=.>r>�>�>�>�>?D?q?�?�?�?�?   @ �   0D0t0�0�0�01&1a1�1�1$2Q2t2�2�2�2!3A3q3�3�3�34!4D4�4�4�4�4$5T5t5�5�56A6a6�6�6�677747]7�7�7848T8t8�8�879�97:q:�:�:�:�:;=;s;�;�;<!<D<�=�=�=>4>k>�>�>�>�>?4?U?t?�?�?�?   P �   010T0t0�0�0141a1�1�1�12242�2�2$3q3�3�3�3�34[4�4�4585S5�5�5�5�5�5666f6�6�6�6�6�6/7C7X7�7�7�7�7898V8k8�8?9�9�9�9P:G<->C>�>�>?P?h? ` �   �0�0�0�011D1d1�1�1�1�1212R2t2�2�2�2U3{3�3d4�4�4Q5d5�5�5�5�56$6A6d6�6�6�6�6717T7t7�7�7D8�8�8�8919Q9t9�9�94:t:�:�:�:;4;T;t;�;�;�;<4<T<�<�<�<�<!=D=q=�=�=�=>A>d>�>�>�>?�?�?   p    u0�0�01�1�1$2�2�2�233-3Q3�3�5K6�6�67K7�7�7�7�7�7�788&898K8]8o8x8�8�8�8�8�89$969T9b9o9�9�9�9�9�9�9�9:#:@:X:r:�:�:�:�:�:�:;;6;H;[;�;�;�;�;�;�;�;�;<%<A<S<p<�<�<�<�<�<�<==5=L=f=x=�=�=�=�=�=�=>=>d>r>>�>�>�>�>�>�>?!?3?P?h?�?�?�?�?�?�?�?   � �   0,0F0X0j0r0�0�0�0�0�01191Z1r1�1�1�12r2z2�2�2�2�2�2�23
33o3�3�3�3�3�4�4�415t5�5�5�5�56646Q6d6�6�6�647"8)80878>8E8L8S8�8�8�8�9	:�:�:�:;/;Q;�;�;<�<�<b=h=�=�=�=�=�=>?>R>l>�>�>�>�>�>�>   �    �7�7�8Q:�:Y;�;�; � L   �45-5e5�5�556u6�6�6"7U7�7�78E8�8�8929b9�9�9:E:�:�:%;e;�;�;%<�<   � �   .1�1�1�1�1�13M3�4�4�45!545d5�5�5�5�5646d6�6�6�6747T7�7�7�7$888G8�8�8�89!9D9d9�9�9�9:!:4:d:�:�:�:<<-<P<>A>d>�>?4?   � �   �0�0�0�0�0 1
1181U1�1�1�1222(212�2�2�2�2�2�2,3S3\3u3�3�3�3�3�364C4M4R4�4�4L5U5�6�6�67%7B7S7]7z7�7�7�78(8i8�8�8�8�8 999%9+969;9&:�:�:�:e=�=�=�=f>n>�>�>�> � (  �0�1�1�1�1�1�1�1�1�12	22222"2(2,22262O2b2�2�2G3a3j3r3�3�3�3w4�4�4�4�45(5/575<5@5D5m5�5�5�5�5�5�5�5�5�5�56$6(6,606�6�6�6�6�6�6�6�67M7T7X7\7`7d7h7l7p7�7�7�7�7�7J88�8�8�8�8�8�8�89!9(9,9094989<9@9D9�9�9�9�9�9::,:3:8:<:@:a:�:�:�:�:�:�:�:�:�:�:*;0;4;8;<;�;�;G<[<�<==2=O=\=�=C?U?   � x   '010>0Y0`0x0�0�0�01W1]1n1�1�1�12!2�2�2�23%3�3�3�3�4�5�5�5�5G6�6�6�7=9�:�;;=E=�=;>@>J>~>�>�>�>�>�>?;?W?o?�?�? � �   T0f0�0�0�01$1<2G2�2�2333q3{3�3�34B4M4_4s4�4�4�4�4�4�4�45�5b6�67�7`8h8�8�8T9`9�9�9W:c:�:�:;�;�=\>n>x>�>�>�>�>�>???S?\?h?�?�?�?�?�?   t   0�0�0�0�1�1�12W23F3�3�3,4t4 55(5d5�5�5�5�5�5�5�5�5�6*7{7�7�7�788p8�8�8�8<9�9�:m;P=�=�=>>o>�>?O?W?    4   �0%191i1s11�1�1v2n3�34q6~6�6Y78x9�9];�<�?   L  0(0&23%303<3Q3X3l3s3�3�3�3�3�3�3�3�3444$43494B4N4\4b4n4t4�4�4�4�4�4�4�4�45+5k5q5�5�5�5�5�5u6�6�6�6�6.7>7D7P7V7f7l7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78888$8*8.84898?8D8S8i8t8y8�8�8�8�8�8�8�8�8�8�8	9%9q9|9�9�9::$:*:0:6:=:D:K:R:Y:`:g:o:w::�:�:�:�:�:�:�:�:�:�:�:�:�:;;;5;:;z<�<�<A>R>�>�>�>�>�>�>�>??&?0?C?g?�?�?�?   0 L   V0s0�0'1F1�1�1�1�1222.2G2c2l2r2{2�2�2�2�2�2%3A3d3w3�4z58s8�8>�> @   d0�0�0�0�0�0�0?1G1T1�1�1!2*2E2Q2]2i2�2�2�2�2�2�2�2�2333"3.3:3C3L3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3F4�45�6777!7-747=7P7Z7f7o7w7�7�7�7�7�7�7�7�7�788,8@8F8O8b8�89;9I9N9�;�;�;�;�;�;�;�;�;<<$<*<0<5<><[<a<l<q<y<<�<�<�<�<�<�<�<�<�<�<�<===)=�=   P �   *161i1�1�12�3�3�3	4&4�4\5d5|5�5�5�566,696E6U6\6k6w6�6�6�6�6�6�67@7O7X7|7�7p8�8�8�899L9�9�9�9�9:6:w:�:�:;;5;S;u;�<�<=m=�=�>�>�?�?   ` T   0�1�2O3�3�3�3�3�4�4�4o5�5�5�56�6�6�7Q8�9E:R:r:�:�:�:�;c<�=>A>K>c>�>�>�>   p    ,0�0�0�0�7   � �   2&2E2N2{2�2�2�2�2�2-353H3S3X3h3r3y3�3�3�3�3�3�3�3�34A4N4x4}4�4�4�475D5L5[5�5�5�5�5666�7�7�7�7�7�7g8m8�8�8�8�8�8�8�8K9^9�9�9�9�9�9�9:�:�:�:�:�;�;�;�;�;�;�;<<-<d<|<�<�<�<�<�<=	=1=V={=�=�=�=�=>>�>�?�?�?   � T   )0<0W0�3�46K6p6S8O:S:W:[:_:c:g:k:{:�:�;�;�; <8<{<�<�<�<l=>>>/>?>K>I?�?   � 8   X0�01^1f1u1}1�129Y:t:�:f;p;�;�;=,=}=!>+>M>? � �   0,0=0E0U0f0u0�0�0�01�1�1)333K3R3\3d3q3x3�3A4�4 5|5�5�5�5�5>6q6�677k7q7�7�7�7�7�7E8�8�8�8�8�8(969}9�9�9�9�9�9�9�9S:\:b:   � l   �0�01/1A1z1�2�2�2�2-3?3Q3c3u3�3�3�3�5606V8l8}8�8�8�8�8�8m9�9:):y:�:K<�<C=L=�=�=�=%>k>t>�>�>�> ?/? �    a4   � �   �5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�566666i6)8`88�8�8999D9z9�9�9�9�9�9 ::a:m:y;<m<y<�<==�>�>�?   � X   �1�5@7[7q7�7�7�79s9�9	:W:h<z<�<�<�<�<�<*=3=H=x=(>->?>]>q>w>�>??4?A?F?T?�?�?     �   {132=2�2 3w3�3\4f45A5u5�56�6�6�6707�7+8F8T8\8i8�8�8�8�8�8�8�8�8�8�9:C:V:g:�:�:�:�:;h;y;�;�;+<6<d<r<{<�<�</=<=d=�=�=�=�>�?�?�?�?�?�?�?�?�?�?�?    `   000!0+090y0�0�0�0�0�0$1/1Z2x2�2�233*323?3F3 44�4�5�68�:y;�;�;<%<8<J<�<�<�?�?�?     P   0-080O0t0�0@1i2e3A475?5�5�6m7s788+8�8�8�9{:�:6;<�<�<Y=_=o=>&>V>�>   0 4   �1�1555!5%5)5-5155595=5A5N5)6A6P6|6�6 7   @ X   
1�2�2�2�2�2�2�3�3O4V4�4�4,56�679&9U9�9�9�9�:;';=;�;�;<A<}<�<�<=2=�=K>�>�? P 4   q2�3�4�58S8�8�8�8H9�9:y:;2;�;�;Y<>F>�?   ` �   �0+1{1�1�1232Z2�2�263d3�3�3	4D4j4�4�405Z5�5�5�5+6Z6�6�6�67J7�7�7�798�8�8�8,9]9�9�9�9:@:c:�:�:�:;;1;=;G;S;_;i;u;�;�;�;�;�;�;�;�;�;�; p �  `1d1h1l1p1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7�7�7<9@9D9H9L9P9T9X9\9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;H;L;\;`;d; <$<(<,<0<�<�<�<�<�< =   � 8   x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5T6X6\6`6�6�6   � x  x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 8888 8(8080>4>8><>@>D>H>L>P>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�? � D  �1�1H2L2\2`2d2l2�2�2�2�2�2�2�2�2�2�2�233 30343H3L3\3`3h3�3�3�3�3�3�3�3�3�3�3�3 44444$4<4@4X4h4l4t4�4�4�4�4�4�4�4�4�4�4�4�45555 585<5T5X5p5�5�5�5�5�5�5�5�5�5�5�5�5�5�566,606@6D6H6P6h6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67 7$74787<7D7\7l7p7�7�7�7�7�7�7�7�7�7�7�7�78888 8$8,8D8T8X8h8l8p8t8|8�8�8�8�8�8�8�8�8�8�8�8�8 999$9(9@9P9T9h9l9|9�9�9�9�9�9�9�9�9�9�9�9�9�9:::,:0:8:P:`:d:t:x:|:�:�:�:�:�:�:�:�:�:�:�: ;; ;0;4;D;H;P;h;x;|;�;�;�;�;�;�;�;�;�;�;�; <<<$<(<8<<<@<H<`<p<t<�<�<�<�<�<�<�<�<�<�<�<�<=== =0=4=8=@=X=h=l=|=�=�=�=�=<?D?P?p?x?�?�?�?�?�?�?�?�?�? � 8   00040<0D0L0T0\0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01111$101T1t1|1�1�1�1�1�1�1�1�1�1�1�1�1 22,242@2`2h2t2�2�2�2�2�2�2�23303<3`3�3�3�3�3�3�3�3�3�3�3�3�3�3�3444$4,444<4D4P4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�45555$5,545<5D5L5T5\5d5l5t5|5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�78888$8,848<8D8L8T8\8d8l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89999(9H9P9X9`9h9p9x9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 ::::<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<= =@=H=T=t=|=�=�=�=�=�=�=�=�=�=>>0>8>@>H>P>X>`>h>t>�>�>�>�>�>�>�>�>�>�>�>??? ?(?0?8?@?H?P?\?|?�?�?�?�?�?�?�?�?�?�?�?�?   � D  0$0,040<0H0h0p0x0�0�0�0�0�0�0�0�0�0�0�0�01 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2L2p2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 3333 3(30383@3H3P3X3`3h3t3�3�3�3�3�3�3�3�3�3�3�3�3�3�34444$4,444<4D4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4555$5,5@5H5T5t5�5�5�5�5�56$646H6X6l6t6�6�6�6�6�6�6 77<7D7L7T7\7h7�7�7�7�7�7�7�7�7�78848<8D8P8p8|8�8�8�8�8�8�8�8�8�8�8 9 9(90949<9P9X9`9h9t9�9�9�9�9�9�9�9::: :@:D:H:P:d:l:�:�:�:�:�:�:�:;$;P;X;|;�;�;�;�;�;�;�;<,<4<@<h<|<�<�<�<�<�<�<�<=$=D=P=x=�=�=�=�=�=�=�= >> >P>\>|>�>�>�>�>�>�>??$?<?t?�?�?�?�?�?�? �    000<0P0h0�0�0�0�0�0�0�0�0�01$101P1X1d1�1�1�1�1�1�1�122$2D2L2T2`2�2�2�2�2�2�2�2 3 3@3L3h3�3�3�3�344(4H4h4�4�4�4�4�4�4�4555<5H5P5�5�5�5�5�5�5�5�5�5�5�5�5 6 6,6H6T6l6p6�6�6�6�6�67707L7P7p7�7�7�7�7808P8p8�8�8�8�8�899,909P9p9�9�9�9�9�9   �    00 080<0@0\0x0�0�0�0�01L1�1�1�102P2�2�2 3 3@3d3�3�3�3�3�3�34 4$4(4D4`4x4�4�4�4�4�4�4�4�4�4�4�4�4554585<5@5D5H5L5P5T5X5\5`5d5h5p5t5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6 777777$70747`7�;�<==(=8=\=h=l=p=t=x=�=�= ???????? ?$?   l  X0`0343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3~4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�455
555555"5&5*5.52565:5>5B5F5J5N5R5V5Z5^5b5f5j5n5r5v5z5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(686@6D6H6L6P6T6X6\6`6d6p6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7,747<7D7L7T7\7d7l7t7|7`9d9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            