MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       }c�9g�9g�9g��(��;g�0��&g�0���g��v�<g�9g�Yg�0��dg�0��8g�0��8g�Rich9g�                PE  L ΁qP        � !	  �        hR     �                         �                              �Y Q   �Q <                            � �;  ��                            8 @            � \                          .text   ��     �                   `.rdata  �y   �  z   �             @  @.data   �;   `     B             @  �.reloc  ^H   �  J   `             @  B                                                                                                                                                                                                                                                                                                                                                                                                U���}V��H�QV�ҡ�}�H�U�AVR�Ѓ���^]� U���}V��H�QV�ҡ�}�U�H�E�IRj�PV�у���^]� ���������̡�}�P�BQ��Y�U��j�h��d�    P��VW�Pg3�P�E�d�    �E�    ��}�P�E���   P�EP�E�P�ҋ���}�H�u�QV�E�   �ҡ�}�H�QVW�ҡ�}�H�A�U�R�E�   �E� �Ѓ��ƋM�d�    Y_^��]� ���������U��W�}��xS�]V�u����u��y�^[_]� ���������U��j�h�d�    PQV�Pg3�P�E�d�    ��u��e �N�E�    ����]` �N$�E��� �ƋM�d�    Y^��]����������������U��j�h!�d�    PQV�Pg3�P�E�d�    ��u�����N$�E�   �2� �N�E� �F` ���E������d �M�d�    Y^��]���������U���T  �Pg3ŉE�Wj j�_ ����u_�M�3��# ��]�V������PWǅ����(  �X_ ����   ������Qj�H_ �����   ������RPǅ����$  �_ ���}   ������P������h  Q�R& ������h  R��% ���������P�I �@��u�+�$    ��/t��t������H��\uꍴ����V�% h�V�R ����u.������PW�^ ���8���W� �^3�_�M�3��" ��]ËM�^3͸   _�x" ��]���������j j j�� �����U��j�h��d�    P��`SVW�Pg3�P�E�d�    ��E�P�M�Q3ۋ��E�   �]��;n 9]��2  �M��Z� ��}�B�P�M�Q�]��҃��E�Pj�M܍~Q���E��Z���P�M��E��� �U�R�M��E���� �M��E���� ��}�H�A�U�R�E��Ћ�}�Q�J�E�P�]��у�h���M���� �U�R�M��E��� �M��]��� �E�SP�r� �����X  ��}�Q�J�E�P�ы�}�B�PSj��M�h��Q�ҍE�P�E��� ��}�Q�J�E�P�]��у�S����d ��}�B�P�M�Q�ҡ�}�H�ASj��U�hx�R�ЍM�jQ�E��$ ��}���B�P�M�Q�E�]��҃� S8]���   hh��M������E�P�E��A ��}�Q�J�E�P�]����� h�h�   h ~h�   �E���� ���E��E�;�t	��覟  �3��U�WR�Ȉ]��s�  h�  ����c �S�E�P���E�   �]��O� �M��E������ � �M�d�    Y_^[��]� ������������U���SVW��j�~W�E�3�P�E�   �]��:� jW�M�Q���E�   �]��"� jW�U�R���E�   �]��m jW�E�P���E�   �]��"m jW�M�Q���E�   �]��
m jW�U�R���E�   �]���l jW�E�P���E�   �]���l jW�M�Q���E�   �]���l j
W�U�R���E�
   �]��
m j	�E�	   �]�W�E�P���l jW�M�Q���E�   �]��zl jW�U�R���E�   �]��bl jW�E�P���E�   �]��� jW�M�Q���E�   �]��2l _^[��]������������U��j�h�d�    P���   SVW�Pg3�P�E�d�    ����� ���  h���M��� ��l���3�P�]���� �M�QP�U�R�E��� ���~$P���E��D� �M��E��� ��l����]���� �M��E�������� �^@�C� �E�SW�E�   �� �����Q  �E�P���|� P�M��E��/� jj�M�Q�M�htaoc�E��6� ���M��E��E��� ��}�B�P�M�Q�E��҃�8]�t'�E�P�E�������� ��3��M�d�    Y_^[��]�Sh���M��!�����}�Q�R8�E�P�~j���E��ҡ�}�H�A�U�R�E��Ѓ�h���M��/� h����l����E��� ��4���j	Q�E��y� ��l���RP��P���P�E�	�� �M�QP�U�R�E�
��� �� ��P����E�荿 ��4����E��~� ��l����E��o� �M��E��c� �E�jP�8� ���M���t8Q�M��� ��}�RP�B8j���E��Ћ�}�Q�J�E�P�E����jSh�������P�E��	 ��}�B�P�M�Q�E��҃�Sh���M��������}�P�R8�E�Pj���E��ҡ�}�H�A�U�R�E��Ћ�}�Q�B4��Sj���Ћ�}�Q�B0jj���Ћ�}�Q�B0jj���Ћ�}�Q�B0Sj���Ћ�}�Q�B0Sj���Ћ�}�Q�B0jj���Ћ�}�Q�B4Sj
���Ћ�}�Q�B0jj	���Ћ�}�Q�B0jj���Ћ�}�Q�B0Sj����Sh���M��������}�Q�E��E�P�R8j���ҡ�}�H�A�U�R�E��Ћ�}�Q�B0��Sj���ЋM�W�z� �M��2� �M��E��v� �M�Q�N$�*� P�M��E��ݼ �M�jj�U�Rhtaoc�E���� ���M��E��E��2� ��}�H�A�U�R�E��Ѓ�8]�t'�M�Q�E������u� ��3��M�d�    Y_^[��]ËM�j�~W�P� �M��� ��}�E�   �]�B�P�M�Q�҃��E�Pj�M�Q���E������SSP�U�R���E��c ��}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��ы�}�E�   �]�B�P�M�Q�҃��E�Pj�M�Q���E��s���SSP�U�R���E��b ��}�H�A�U��E�R�Ћ�}�Q�J�E�P�E��ы�}��h���h  �Sjh���h  ��E�   �]�B���   Sj����P�E�P���p^ ��}S�E�   �]�Q���   Sj����P�M�Q��裧 ��}S�E�   �]�B���   Sj����P�E�P���v� ��}S�E�   �]�Q���   Sj����P�M�Q���I� ��}SS�E�   �]�Bj���   ����P�E�P���� ��}S�E�   �]�Q���   Sj����P�M�Q���� ��}h���h  �Sjh���h  ��E�
   �]�B���   Sj
����P�E�P���L] ��}S�E�	   �]�Q���   Sj	����P�M�Q���� ��}S�E�   �]�B���   Sj����P�E�P���R� ��}S�E�   �]�QSj�ϋ��   ��P�M�Q���%� ��}�E�   �]�B�P�M�Q�҃��E�Pj�M�Q���E�����SSP�U�R���E��?` ��}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��ы�}��S�E�   �]�B���   Sj����P�E�P��脥 h�  ����Y �M�Q�E������� ���   �M�d�    Y_^[��]���������������U��j�h��d�    P��0VW�Pg3�P�E�d�    ���@ ��   �H� �E��E�P�O$�E�    蒹 P�M��E��E� jj�M�Q�M�htaoc�E��L� �Mċ��E�螸 ��}�B�P�M�Q�E� �҃���t���z����M���W�^� �M��� �E�P�E�������� ���M�d�    Y_^��]���U��j�hL�d�    P��   SVW�Pg3�P�E�d�    ��3ۉ]��F@   �����E����   ����   ���"  ��}�H�A�U�R�Ћ�}�Q�JSj��E�hh�P�эU�R�E�   �9 ��}�H�A�U�R�E��������� h�h�   h ~h�   ����� ��,�E�E�   ;�t	��虓  �3���VW���E������b�  �{  �MQ�U�R���E�   �]��` 9]�Y  h�  ���W �H  �%� h�h�   h ~j$���]� ��;�t�@   ��X�X�X�X�3���VW���E������H  ��}�H�A�U�R�Ѓ��M�Qj�Uؿ   R�Ή}��������}�H�A�U�R�E��Ћ�}�Q���   ��Sj���Ѕ�t2Sh���M��=�����}�Q�Rx�E�P�M��E��}����E��u�]�E��E�   t��}�H�A�U�R�Ѓ�8]�  ���������   ��}�Q�BdW�M��Ћ�}�Q�����   h��h�   V�Ћ�}�Q��j���BhVW�M���j<��L���SQ�� ����L���RǅL���<   ��P�����T���ǅX���4���\�����d���ǅh���   ��l����T���ufSh��M��&����E�P�E��� ��}�Q�J�E�P�E����0Sh��M�������U�R�E��� ��}�H�A�U�R�E��Ѓ���}�Q�J�E�P�E������у��   �M�d�    Y_^[��]� ���������V��V�� ���    ^�������������U��V�������Et	V�� ����^]� �������������������P�P�����U������P�M�P��P(�P �P�P@�P8�P0�PX�PP�XH���Q�P�Q�P�Q�P�Q�P�I�H�M��P�Q�P�Q�P �Q�P$�Q�P(�I�H,�M��P0�Q�P4�Q�P8�Q�P<�Q�P@�I�HD�M��PH�Q�PL�Q�PP�Q�PT�Q�PX�I�H\]� �����������U��M�U�A�
�E��B�I0���B�IH����A �
�A�A8�J���AP�J���X�A(�
�A�A@�J���AX�J���X�A�J�B �I0���B(�IH���X�A8�J �A �J���AP�J(���X �A@�J �A(�J���AX�J(���X(�A�J0�A0�J8���AH�J@���X0�A8�J8�A �J0���AP�J@���X8�A@�J8�A(�J0���AX�J@���X@�A�JH�BP�I0���BX�IH���XH�BP�I8�BH�I ���AP�JX���XP�A@�JP�BH�I(���AX�JX���XX]�������������������U���}�UV��H�AVR�Ѓ���^]� ��������������U��j�h��d�    P��VW�Pg3�P�E�d�    �U�E�    ��}�H�I(R�E�P�ы���}�B�u�HV�E�   �ы�}�B�HVW�ы�}�B�P�M�Q�E�   �E� �҃��ƋM�d�    Y_^��]����������������U��j�h��d�    P��VW�Pg3�P�E�d�    �U �E�E�    ��}�H�ER�UP�ERP�A$���U��$R�Ћ���}�Q�u�BV�E�   �Ћ�}�Q�BVW�Ћ�}�Q�J�E�P�E�   �E� �у�,�ƋM�d�    Y_^��]����������̡�}���   �Q��Y���������������U��j�h��d�    P��$SVW�Pg3�P�E�d�    3ۉ]Љ]؋E�M�Q�M�]��E��]�]��� �}S�U�R�E�P���E���& �M���]��A ;�tz��}���   �JX�E�P�ы���;�t\��}���   �PT���ҋ�}�Q|�M�RQPV�ҋ��}���   ��U�R�E������Ѓ��ƋM�d�    Y_^[��]� ��}���   �
�E�P�E������у�3��M�d�    Y_^[��]� ���������������U��j�h�d�    P��(SVW�Pg3�P�E�d�    3ۉ]��]̉]ԋE�M�Q�   �M�}��E܉]��]�� �MS�U�R�E�P�E��% �M���E��
 ;�t\��}���   �JH�E�P�ы�}�u���B�HV�ы�}�B�HVW�ы�}���   ��M�Q�E�   �]��҃��C��}�H�u�QV�ҡ�}�H�QSj�h��V�ҡ�}���   ��U�R�}��]��Ѓ��ƋM�d�    Y_^[��]� �U��j�h/�d�    P��$SV�Pg3�P�E�d�    3ۉ]Љ]؋E�M�Q�M�]��E��]�]�� �MS�U�R�E�P�E��q$ �M���]��� ;�tJ��}���   �J8�E�P�ы�}�����   ��M�Q�E������҃��ƋM�d�    Y^[��]� ��}���   ��U�R�E������Ѓ�3��M�d�    Y^[��]� ����U��j�hk�d�    P��(SV�Pg3�P�E�d�    3��u��ủuԋE�M�Q�M�u��E܉u��u�� �MV�U�R�E�   P�]��]��w# ��t��}���   �J�E�P�у���u2ۍM�u��� ��t7��}���   �P<�M�Q���]��}���   ��U�R�E������Ѓ����}���   �
�E�P�E������у��E�M�d�    Y^[��]� �����������U��j�h��d�    P��$SV�Pg3�P�E�d�    3ۉ]Љ]؋E�M�Q�M�]��E��]�]�� �MS�U�R�E�P�E��q" �M���]��� ;�tZ��}���   �J@�E�P�ыu��H��P�N�H�V�P�@�N��}�V���   �
�F�E�P�E������у��+���}�u�V���   �V���M�Q�E������҃��ƋM�d�    Y^[��]� ������U��j�hڳd�    P��(SV�Pg3�P�E�d�    3ۉ]��]̉]ԋE�M�Q�M��E�   �E܉]��]��o �MS�U�R�E�P�E��Z! �M���E��� ;�tC��}���   �JL�E�P�ыu��P���� ��}���   ��M�Q�E�   �]����(�uS���j� ��}���   ��U�R�E�   �]��Ћƃ��M�d�    Y^[��]� �����U��j�h��d�    PQSVW�Pg3�P�E�d�    ��}�P�Bd3�j�M�}��Ћ�}�Q�����   hH�Fh�  V�Ћ�}��j�E��QVP�Bh�M��N;�~�]��M��R��葲 G;�|�E�P��� ��}�Q�J�EP�E������у��M�d�    Y_^[��]� ���U��j�h �d�    P��SVW�Pg3�P�E�d�    ��}�H�A�U�R�Ћ�}�Q�J3�Wj��E�h��P�у���}�B�Pdj�M��}��ҋ��}�H���   hH�Fh�  V�ҋ�}��j�E��QVP�Bh�M���N;�~�]��M��R��葱 G;�|�E�P��� ��}�Q�J�E�P�E������у��M�d�    Y_^[��]� ���U��Q�ESVW���   3�3�3�3ۃ��M�|#�@|�O���A�	�d$ p����u�E�M�;�}�@|��_�^�[��]� �����U��j�h��d�    P��   SV�Pg3�P�E�d�    3ۉ]��}�H�u�QV�]��ҡ�}�H�QSj�h8�V�҃��E�]��E�   ��
�j  �$��4 Sh4��M��)����E�P���E�   �[  ��}�Q�J�E�P�]����&  Sh0��M�������U�R���E�   �m[  �U���  Sh(��M�������M�Q���E�   �E[  ��}�B�P�M�Q�]�����  Sh$���p���������p���P���E�   �[  ��}�Q�J��p���P�]����  Sh ��M��J����U�R���E�   ��Z  �U��H  Sh���P���������P���Q���E�   �Z  ��}�B�P��P���Q�]����  Sh��M�������E�P���E�   �]Z  ��}�Q�J�E�P�]�����   Sh��M������U�R���E�   �#Z  �U��   Sh��M��}����M�Q���E�	   ��Y  ��}�B�P�M�Q�]����}Sh����`����C�����`���P���E�
   �Y  ��}�Q�J��`���P�]����=Sh����@���������@���R���E�   �~Y  ��@�����}�H�AR�]��Ѓ���}�Q�J�E�P�ы�}�B�PSj��M�h��Q�҃���}�P�B<���E�   �Ћ�}�Q�RLj�j��M�QP���ҡ�}�H�A�U�R�]��Ѓ��ƋM�d�    Y^[��]� ���1 32 [2 �2 �2  3 C3 }3 �3 �3 4 ������������U��j�h9�d�    PQSVW�Pg3�P�E�d�    ���}�3��   �G�7�w�w�w�w�_�u��C�3�s�s�s�s�G@�w0�w4�wD�w<�w8�GX�wH�wL�w\�wT�wP�Gp�w`�wd�wt�wl�wh���   �wx�w|���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   �E�97t	W�� ���7�w�w�w�w93t	S�q� ���G0�3�s�s�s�s90t	P�S� ���GH�w0�w4�wD�w<�w890t	P�4� ���G`�wH�wL�w\�wT�wP90t	P�� ���Gx�w`�wd�wt�wl�wh90t	P��� �����   �wx�w|���   ���   ���   90t	P�˿ �����   ���   ���   ���   ���   ���   90t	P蚿 �����   ���   ���   ���   ���   ���   �ǋM�d�    Y_^[��]����������������U��j�h��d�    PQSVW�Pg3�P�E�d�    ��u��E�   ��� ���   3��E�9t	W�� ����_�_�_�_���   �E�9t	W�޾ ����_�_�_�_�~x�E�9t	W輾 ����_�_�_�_�~`�E�9t	W蚾 ����_�_�_�_�~H�E�9t	W�x� ����_�_�_�_�~0�E�9t	W�V� ����_�_�_�_�~�]�9t	W�5� ����_�_�_�_�E�����9t	V�� ����^�^�^�^�M�d�    Y_^[��]�U��j�h��d�    P��(  SVW�Pg3�P�E�d�    ���}��}�H�A�U�R�Ћ�}�Q�Jj j��E�hX�P�ы�}�B�P��|���Q�E�    �ҡ�}�H�Aj j���|���hL�R�ЋMQ�����R�E������P��|���P��<���Q�E��[  �U�RP�E�P�E��[  ��H��}�Q�J��<���P�E��ы�}�B�P�����Q�E��ҡ�}�H�A��|���R�E��Ћ�}�Q�J�E�P�E��ы]��}�B�H��S����e�V�ы�}�B�P�M�VQ�҃��������u�F�E�    ���k  3���}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�ы�}�B�P�M�Q�E�	�ҡ�}�H�Aj j��U�hH�R�Ћ�}�Q�J��\���P�E�
�ы�}�B�Pj j���\���hH�Q�ҡ�}�H�A�U�R�E��Ћ�}�Q�J��@j j��E�hD�P�у��F�D8j0j j�j ���U��$�E�R��������؋F�D8j0j j�j ����L����$P�E��������E�F�8j0j j�j ����l����$Q�E��s���P�U�R��,���P�E��Y  ��\���QP������R�E��vY  �MQP������R�E��aY  ��@�M�QP�����R�E��IY  SP������P�E��7Y  �M�QP������R�E��"Y  ��}�Q�R�M�QP�E��ҡ�}�H�A������R�E��Ћ�}�Q�J������P�E��ы�}�B�P�����Q�E��ҡ�}�H�A������R�E��Ћ�}�Q�J������P�E��ы�}�B�P��,�����@Q�E��ҡ�}�H�A��l���R�E��Ћ�}�Q�J��L���P�E��ы�}�B�P�M�Q�E��ҡ�}�H�A�U�R�E����E�
��}�Q�J��\���P�ы�}�B�P�M�Q�E�	�ҡ�}�H�A�U�R�E��ЋM��}�B�� Q�H���܉eS�ы�}�B�P�M�SQ�ҋM�������E�@��;F�E�������}�]��}�H�A�U�R�Ћ�}�Q�Jj j��E�hX�P�ы�}�B�P�M�Q�E��ҡ�}�H�Aj j��U�h<�R�ЋMQ��l���R�E��/���P�E�P��L���Q�E���V  �U�RP�E�P�E���V  ��H��}�Q�R�M�QP�E��ҡ�}�H�A�U�R�E��Ћ�}�Q�J��L���P�E��ы�}�E��B�P��l���Q�ҡ�}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��ы�}�B�H��S����eV�ы�}�B�P�M�VQ�҃����D���S��������}�H�A�U�R�E������Ѓ��M�d�    Y_^[��]� �������������U��j�h\�d�    P��  SVW�Pg3�P�E�d�    ���}��}�H�A������R�Ћ�}�Q�Jj j�������ht�P�ы�}�B�P�����Q�E�    �ҡ�}�H�Aj j������hL�R�Ћu�F,P������Q�E��N���P�����R��(���P�E��U  ������QP�U�R�E��U  ��H��}�H�A��(���R�E��Ћ�}�Q�J������P�E��ы�}�B�P������E�Q�ҡ�}�H�A������R�E��ЋM��}�B��Q�H���܉eS�ы�}�B�P�M�SQ�҃�������3�9]�]�  ��}�H�A������R�Ћ�}�Q�Jj j�������h��P�ы�}�B�P��x���Q�E�	�ҡ�}�H�Aj j���x���hH�R�Ћ�}�Q�J������P�E�
�ы�}�B�Pj j�������hH�Q�ҡ�}�H�A������R�E��Ћ�}�Q�J��@j j�������hp�P�у��Fj0�<[�j �j�j ��E����@��(����$R�������E���F�d8j0j �jj ��������$P�E���������E�F�8j0j j�j ���������$Q�E�����P������R��x���P�E���R  ������QP��H���R�E��R  �M�QP��H���R�E��R  ��@��x���QP��h���R�E��R  �M�QP��X���R�E��yR  �E�������QP��x���R�aR  ��}�Q�R�M�QP�E��ҡ�}�H�A��x���R�E��Ћ�}�Q�J��X���P�E��ы�}�B�P��h���Q�E��ҡ�}�H�A��H���R�E��Ћ�}�Q�J��H���P�E��ы�}�B�P��x�����@Q�E��ҡ�}�H�A������R�E��Ћ�}�Q�J�����P�E��ы�}�B�P��(���Q�E��ҡ�}�E��H�A������R�Ћ�}�Q�J������P�E�
�ы�}�B�P��x���Q�E�	�ҡ�}�H�A������R�E��ЋM��}�� Q�J�Q���ĉe�P�E��ҡ�}�H�U��IR�E�P�ыM���������}�B�P������Q�ҡ�}�H�Aj j�������h��R�Ћ�}�Q�J�E�P�E��ы�}�B�Pj j��M�hH�Q�ҡ�}�H�A������R�E��Ћ�}�Q�Jj j�������hH�P�ы�}�B�P��X���Q�E��ҡ�}�H�A��@j j���X���hp�R�Ѓ��N�D(j0j j�Dj ����h����$R�E��������E���F�d j0j j�Dj ���������$Q�E��g������E��V�Dj0j j�|j ���$�E�������P�8���P��X���Q������R�E��PO  ������QP������R�E��8O  �M�QP�����R�E��#O  ��@�M�QP������R�E��O  �M�QP������R�E� ��N  ������QP������R�E�!��N  ��}�Q�R�M�QP�E�"�ҡ�}�H�A������R�E�!�Ћ�}�Q�J������P�E� �ы�}�B�P������Q�E��ҡ�}�H�A�����R�E��Ћ�}�Q�J������P�E��ы�}�B�P��������@Q�E��ҡ�}�H�A������R�E��Ћ�}�Q�J������P�E��ы�}�B�P��h���Q�E��ҡ�}�H�A��X���R�E��Ћ�}�Q�J������P�E��ы�}�B�P�M�Q�E��ҡ�}�H�A������R�E��ЋM��}�B�� Q�H�����e�W�ы�}�B�P�M�WQ�ҋM���k�����}�H�A��h���R�Ћ�}�Q�Jj j���h���h��P�ы�}�B�P�M�Q�E�#�ҡ�}�H�Aj j��U�hH�R�Ћ�}�Q�J�E�P�E�$�ы�}�B�Pj j��M�hH�Q�ҡ�}�H�A�����R�E�%�Ћ�}�Q�J��@j j������hp�P�у��E�&�Fj0�|[�j �j��D8�j ����x����$R�������E���F�d8j0j �jj ���������$P�E�'��������E��F�8j0j j�j ���������$Q�E�(�����P�����R������P�E�)��K  �M�QP������R�E�*��K  �M�QP�����R�E�+�K  ��@�M�QP��8����E�,R�K  �M�QP��X���R�E�-�K  ��h���QP��h���R�E�.�iK  ��}�Q�R�M�QP�E�/�ҡ�}�H�A��h���R�E�.�Ћ�}�Q�J��X���P�E�-�ы�}�B�P��8���Q�E�,�ҡ�}�H�A�����R�E�+�Ћ�}�Q�J������P�E�*�ы�}�B�P��������@Q�E�)�ҡ�}�H�A������R�E�(�Ћ�}�Q�������E�'P�J�ы�}�B�P��x���Q�E�&�ҡ�}�H�A�����R�E�%�Ћ�}�Q�J�E�P�E�$�ы�}�B�P�M�Q�E�#�ҡ�}�H�A��h���R�E��ЋM��}�B�� Q�H�����e�W�ы�}�B�P�M�WQ�ҋM��������N|�E�<��t  ��}�B�P�M�Q�ҡ�}�H�Aj j��U�h��R�Ћ�}�Q�J�E�P�E�0�ы�}�B�Pj j��M�hH�Q�ҡ�}�H�A��(���R�E�1�Ћ�}�Q�Jj j���(���hH�P�ы�}�B�P��H���Q�E�2�ҡ�}�H�A��@j j���H���hp�R�Ѓ��Fj0�|[	�j �j�j ��E�3���@��8����$Q�������E���F�d8j0j j�j ���������$R�E�4�k������E��F�8j0j j�j ���������$P�E�5�?���P��H���Q������R�E�6�WH  ��(���QP������R�E�7�?H  �M�QP������R�E�8�*H  ��@�M�QP�����R�E�9�H  �M�QP��8���R�E�:��G  �E�;�M�QP��X���R��G  ��}�Q�R�M�QP�E�<�ҡ�}�H�A��X���R�E�;�Ћ�}�Q�J��8���P�E�:�ы�}�B�P�����Q�E�9�ҡ�}�H�A������R�E�8�Ћ�}�Q�J������P�E�7�ы�}�B�P��������@Q�E�6�ҡ�}�H�A������R�E�5�Ћ�}�Q�J������P�E�4�ы�}�B�P��8���Q�E�3�ҡ�}�E�2�H�A��H���R�Ћ�}�Q�J��(���P�E�1�ы�}�B�P�M�Q�E�0�ҡ�}�H�A�U�R�E��ЋM��}�B�� Q�H�����e�W�ы�}�B�P�M�WQ�ҋM���x����E�N|�@;E�E������}��}�B�P�M�Q�ҡ�}�H�Aj j��U�ht�R�Ћ�}�Q�J�E�P�E�=�ы�}�B�Pj j��M�h<�Q�ҋv,������VP�E�>�����P�M�Q������R�E�?�E  �M�QP��8����@R�]��E  ��H��}�Q�R�M�QP�E�A�ҡ�}�H�A��8���R�]��Ћ�}�Q�J������P�E�?���E�>��}�B�P������Q�ҡ�}�H�A�U�R�E�=�Ћ�}�Q�J�E�P�E��ы]��}�B�H��S����eV�ы�}�B�P�M�VQ�҃��������S���������}�H�A�U�R�E������Ѓ��M�d�    Y_^[��]� ���U��j�h��d�    P���   SVW�Pg3�P�E�d�    ���}�HH�U��p  j h�  R�Ћ�}�Q�}��j �E����   j���Ћ�}�Qj �E����   j���Ћ�}�Q�J���E�P�}��у��E�    ���4  �~ �*  ��\���� � ��0���R�E�� � ���)� P��\����E��ي ��0����E�躇 ��}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�у��U�R��\����E��(� ��}�H�A�U�R�E��Ћ�}�Q�J�E�P�ы�}�B�Pj j��M�h��Q�ҡ�}�H�A�U�R�E��Ћ�}�Q�Jj j��E�h��P�у�,�E���0���R��\���譈 �M�Q���E�螇 P�U�R�E�P�E��B  �M�QP�U��R�]��B  ��}�Q�R�M�QP�E�	�ҡ�}�H�A�U�R�]��Ћ�}�Q�J�E�P�E��ы�}�B�P�M�Q�E��҃�,��0����E��P� ��}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��ы]��S���e����}�B�HW�ы�}�B�P�M�WQ�҃��������S���������\����E� �Ӆ ��]��}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�ы�}�B�P�M�Q�E�
�ҡ�}�H�Aj j��U�h��R�Ѓ�(��}���   �M�Bx�E���P�M�Q�U�R�9A  �M�QP�U�R�E��'A  ��}�Q�R�M�QP�E��ҡ�}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��ы�}�B�E�
�MċPQ�ҡ�}�H�A�U�R�E� �Ћ�}�Q�B��0S�����eW�Ћ�}�Q�J�E�WP�у�������S���j����U�}RWS��������}� t�E��MPQWS���s�����}�B�P�M�Q�ҡ�}�H�Aj j��U�h��R�Ћ�}�Q�J�E�P�E��ы�}�B�Pj j��M�hL�Q�ҋEP�M�Q�E�����P�U�R�E�P�E���?  �M�QP�U�R�E���?  ��H��}�Q�R�M�QP�E��ҡ�}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��ы�}�E��B�P�M�Q�ҡ�}�H�A�U�R�E��Ћ�}�Q�J�E�P�E� �ы�}�J�Q��S���ĉeP�E�ҡ�}�H�U�IR�E�P�у���������}�B�P��L���Q�E    �ҡ�}�H�Aj j���L���h��R�Ћ�}�Q�J��x���P�E��ы�}�B�Pj j���x���h��Q�҃�(�} �E��E    �  �}� ��  �~ ��  ���   �M�������   ��}��� ���   �ȋBx�Ћ�}�Q�R��x���QP�ҡ�}�P�Rx����L���P��x����҅��^  ��}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�ы�}�B�P�M�Q�E��ҡ�}�H�Aj j��U�h��R�Ѝ�x���Q�U�R�� ���P�E��=  �M�QP�� ���R�E��n=  ��@��}�Q�R�M�QP�E��ҡ�}�H�A�� ���R�E��Ћ�}�Q�J�� ���P�E��ы�}�B�P�M�Q�E����E���}�H�A�U�R�Ћ�}�Q��S���ĉe�EP�B�Ћ�}�Q�E�RP�M�Q�҃����������}�H�I��L���R��x���P�у���}�B�P�����Q�ҡ�}�H�Aj j������h��R�Ћ�}�Q�R�E�P�����Q�E��ҡ�}�H�A�����R�E��ЋO|�U�� �<� �E    ��  �]�ۍd$ ��}�H�A�U�R�Ћ�}�Q�Jj j��E�hH�P�у���}�B�P<�M��E��ҋ�}�Q�RLj�j��M�QP�M��ҡ�}�H�A�U�R�E��ЋG4��VÍDP��<���Q�������E��}�B�P<�M��E��ҋ�}�Q�M�RLj�j�QP�M��ҡ�}�H�A��<���R�E��Ѓ��}� ��   �\ ��   ��}�Q�J�E�P�ы�}�B�Pj j��M�h��Q�҃���}�P�B<�M��E��Ћ�}�Q�RLj�j��M�QP�M��ҡ�}�H�A�U�R�E��ЋGL�N�ÍDP��h���Q�������E��}�B�P<�M��E��ҋ�}�Q�M�RLj�j�QP�M��ҡ�}�H�A��h���R�E��Ѓ��E�O|�U@��;��E�����]��}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�у���}�B�P<�M��E��ҋ�}�Q�RLj�j��M�QP�M��ҡ�}�H�A�U�R�E��Ћ�}�Q��S���ĉe�EP�B�Ћ�}�Q�E�RP�M�Q�҃��������E�O|��U@;E�E�������}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�ы�}�B�P�M�Q�E��ҡ�}�H�Aj j��U�h<�R�ЋMQ�� ���R�E� ����P�E�P��<���Q�E�!��8  �U�RP��h���P�E�"�8  ��H��}�Q�R�M�QP�E�#�ҡ�}�H�A��h���R�E�"�Ћ�}�Q�J��<���P�E�!�ы�}�E� �B�P�� ���Q�ҡ�}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��ы�}�B�H��S�����eW�ы�}�B�P�M�WQ�҃�������S���������}�H�A��x���R�E��Ћ�}�Q�J��L���P�E� �ы�}�B�P�M�Q�E������҃��M�d�    Y_^[��]� ��������������U��j�hλd�    P��  SVW�Pg3�P�E�d�    ���}�H�A��P���R�E�    �Ћ�}�Q�Jj j���P���hH�P�э�P���R�EP�M�Q�E��7  ��}�B�P��P���Q�E��ҋE�]��$PS�M�Q���������}�B�P�M�Q�ҡ�}�H�Aj j��U�h��R�Ћ�}�Q�J�E�P�E��ы�}�B�Pj j��M�hH�Q�ҡ�}�H�E���`����AR�Ћ�}�Q�Jj j���`���hH�P�у�<�E�j0j jj ����|����$R�E�����������E�j0j jj ���E��$P�E���������E�E�j0j jj ����@����$Q�E�������`���RP������P�E�	�5  �MQP�����R�E�
�5  �M�QP�����R�E��5  ��@�E�WP��$���P�{5  �M�QP������R�E��f5  ������}�P�B<�M��E��Ћ�}�Qj�j�WP�BL�M��Ћ�}�Q�J������P�E��ы�}�B�P��$���Q�E��ҡ�}�H�A�����R�E��Ћ�}�Q�J�����P�E�
�ы�}�B�P������Q�E�	�ҡ�}�H�A��@���R�E��Ћ�}�Q�J�E�P�E��ы�}�E��B�P��|���Q�ҡ�}�H�A��`���R�E��Ћ�}�Q�J�E�P�E��ы�}�B�P�M�Q�E��ҋE��}�Q��,P�B�����eW�Ћ�}�Q�J�E�WP�у��������Uh�  RS����������  h�  P��4���P��������M��E���v ��M��]���v ����p���Q�M�E�蹥 �U�RW��4���QP�E��C� ����p����E��w �M��]��vw ��}�B�P�M�Q�ҡ�}�H�Aj j��U�hH�R�Ћ�}�Q�J�E�P�E��ы�}�B�Pj j��M�h��Q�ҍEP�M�Q�U�R�E���2  �E��M�QP��|���R��2  ��@��}�Q�R�M�QP�E��ҡ�}�H�A��|���R�E��Ћ�}�Q�J�E�P�E��ы�}�B�P�M�Q�E��ҡ�}�H�A�U�R�]��Ћ�}�Q�J�E�P�ы�}�B�Pj j��M�h��Q�҃�,�E�P�M��E���v �M�QP��|���R�E��2  ������}�P�E��MԋB<�Ћ�}�Qj�j�WP�BL�M��Ћ�}�Q�J��|���P�E��ы�}�B�P�M�Q�E��ҡ�}�H�A�U�R�]��ЋM��}�B��Q�H�����eW�ы�}�B�P�M�WQ�҃��������M��E��nu ��4����E��_u ��}�H�A�U�R�E� �Ћ�}�Q�J�EP�E������у��M�d�    Y_^[��]�$ ����������U��j�h��d�    P���   SVW�Pg3�P�E�d�    ��M���s ��}�H�A�U�R�E�    �Ѓ��M�Q�M�   S�U�R�E�����P��D����]��t ��D���P�M��E��tw ��D����]��vt ��}�Q�J�E�P�E��ы�}�B�P�M�Q�E� �ҋM����D���P舡 P�M��E��;w ��D����E� �t ��}�Q�J�E�P�ы�}�B�Pj j��M�h��Q�҃��E��E�P�M��v ��}�Q�J�E�P�E� �у��U�R�M��wt P�E��=� ��}�H�A�U�R�E� �Ѓ��`x �E�h1D4ChCD4C�E����ؼ Pj S�M�Q���yx ��u;�U�R�E��9x ���M��E�    �E������@s 3��M�d�    Y_^[��]� �~ �E    ��  �F�M��}�<��B�P�M�Q�ҡ�}�H�A��p���R�E��Ћ�}�Q�Jj j���p���h��P�ы�}�B�P�M�Q�E�	�ҡ�}�H�Aj j��U�h�R�Ѓ�,��}���   �Bx���E�
��P�M�Q��P���R�].  ��p���QP��4���R�E��E.  ��}�Q�R�M�QP�E��ҡ�}�H�A��4���R�E��Ћ�}�Q�J��P���P�E�
�ы�}�B�P�M�Q�E�	�ҡ�}�H�A��p���R�E��ЋM���}�B��0Q�H���܉e�S�ы�}�B�P�M�SQ�҃���������}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�ы�}�B�@�M�Q�U�R�E��Ћ�}�Q�J�E�P�E��ыU��}�� R���e�܋H�QS�ҡ�}�H�A�U�SR�Ѓ�������h�  W��������tL��}�Q�B���܉e�S�Ћ�}�Q�Bj j�h��S�ЋM��U��h4  h@  WQR���"���h�  W��������tJ��}�H�Q���܉e�S�ҡ�}�H�Qj j�h��S�ҋE��M��h�	  hD  WPQ���������}�B�P��`���Q�ҡ�}�H�Aj j���`���h��R�Ћ�}�Q�R�E�P��`���Q�E��ҡ�}�H�A��`���R�E��ЋM���}�B�� Q�H�����e�W�ы�}�B�P�M�WQ�҃����������}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�ы�}�B�@�M�Q�U�R�E��Ћ�}�Q�E��J�E�P�ыU��}�H�� R�Q�����e�W�ҡ�}�H�A�U�WR�Ѓ����0�����}�Q�J�E�P�ы�}�B�Pj j��M�h��Q�ҡ�}�H�I�U�R�E�P�E��ы�}�B�P�M�Q�E��ҋE���}�Q�� P�B�����e�W�Ћ�}�Q�J�E�WP�у��������U�R���^�����}�H�A�U�R�E��ЋE@��;F�E�=����M��~s �M�Q�E� �!s ���M��E�    �E������(n �   �M�d�    Y_^[��]� ���������������U��j�h��d�    P��  SVW�Pg3�P�E�d�    �ى�����hG  �c� �K 3����������;���  �������l ��}�H�A�U�R�}��Ѓ��u�M�Qj�U�R���E�豤��P��t����E���l ��t���P�������E��;p ��t����E��<m ��}�Q�J�E�P�E��ы�}�B�P�M�Q�E� �ҋM����t���P�N� P�������E���o ��t����E� ��l ��}�Q�J�� ���P�ы�}�B�PWj��� ���h`�Q�҃��E��� ���P�������Do ��}�Q�J�� ���P�E� �у���8����}k ��}�B�P�M�Q�E��҃��E�Pj�M�Q���E�����P��t����E��k ��t���R��8����E�	�	o ��t����E��
l ��}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��у�hT���t����k ��t���R��8����E�
��n ��t����E��k �������j ��}�H�A�U��E�R�Ѓ��M�Qj�U�R���E�询��P��t����E���j ��t���P�������E��9n ��t����E��:k ��}�Q�J�E�P�E��ы�}�B�P�M�Q�E��҃�hH���t����;j ��t���P�������E���m ��t����E���j �M�Q�������k P�E��M� ��}�B�P�M�Q�E��҃��E�P��8����Uk P�E��� ��}�Q�E��E�P�J�у��U�R�������#k P�E��� ��}�H�A�U�R�E�����ݕx������U���x����@�Q�]��U�R��T����U�P�荍l����U�QݝT����������U�ݕ\���ݕd���ݕl���ݕt���ݝ|���蚵����}���   ���   �щE�MWP�E��u� ��}���   �M䋐�   �҅���  �an �E�h1D4ChCD4C�E��E��ز �M�PWj������P�un ��ux�M�Q�E��4n ��}�}����   ���   �M�Q�E��҃��}䍍�����E�� i ��8����E� �i �������E�������h 3��M�d�    Y_^[��]� Wh���M��˟���E�P�M�Q�������E��i ���ԉe̍M�QPR�E��$  ����賾����}�B�P�M�Q�E��ҡ�}�H�A�U�R�E��Ѓ�Wh���M��W����M�Q�U�R��8����E��i ���̉e̍U�RPQ�E��)$  �����?�����}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��у�Wh���M������U��}R�P���   Wj���E���P�M�Q���
������ԉe̍M�QPR�E��#  ����蹽����}�B�P�M�Q�E��ҡ�}�H�A�U�R�E��Ћ�}�Q���   ��Wj����;�t�M�Q���̉e�Wh0��:������S�����}�B���   Wj����;�t�E�P���̉e�Wh �������������}�Q���   Wj����P�M�Q���)���P�E��o� ��}�B�P�M�Q�E��ҋM�����k Wh��M�蠝��Wh��M��E�莝��������P�������E��Hg P�M�Q������R�E��c"  �M�QP������R�E��N"  P�E� �� ��}�H�A������R�E��Ћ�}�Q�J������P�E��ы�}�B�������E�Q�P�ҡ�}�H�A�U�R�E��Ћ�}�Q�J�E�P�E��у�0�j �E�h1D4ChCD4C�E�!�E��� �M�PWj������R�j ��u4�E�P�E��zj �M�Q�}��E��jj ���M�}��E��x  �D�����}�B�P�� ���Q�҃�Wh���M��E�"�9�����}�H�I�� ���R�E�P�E�#�ы�}�B�P�M�Q�E�"�ҋE��P���� ����̉e�R輛���������   �E���|�����x���Pǅx����  �}��}��}��� ��Wh���M�觛��Wh���M��E�$蕛����x���Q������h��R�E�%�� P�E�P������Q�E�&�d   �E�'�U�RP������P�O   ��$P�� ����E�(�,�����}�Q�J������P�E�'�ы�}�B�P������Q�E�&�ҡ�}�H�A������R�E�%�Ћ�}�Q�J�E�P�E�$�ы�}�B�P�M�Q�E�"�ҋE��P���� ����̉e�R�{������Ĺ��Wh���M�薚��Wh���M��E�)脚����}� P������Q�E�*茱��P�U��E�+R������P�W  �M�QP������R�E�,�B  �� P�� ����E�-������}�H�A������R�E�,�Ћ�}�Q�J������P�E�+�ы�}�B�P������Q�E�*�ҡ�}�H�A�U�R�E�)�Ћ�}�Q�J�E�P�E�"�ыU��R���� ����̉e�P�o�����踸���M�Q���}�����}�B���   Wj���ҋM�{�{�E���}���   ���   �}��Ѕ���  設 ��}���   �E��M䋒�   P�ҋ�}���   �EЋȋB��=�  �#  ��}�Q�J������P�ы�}�B�PWj�������h��Q�҃���}���   �uЋBx���E�.��P������Q��t���R�  P�E�/�0� ��}�H�A��t���R�E�.�Ћ�}�Q�J������P�E�"�у���t����Q�����}�B�P������Q�E�0�ҡ�}�H�AWj�������h��R�Ѓ���}���   �Bx���E�1��P������Q��\���R��  P�E�2蔫 ��}�H�A��\���R�E�1�Ћ�}�Q�J������P�E�0�у�9}���  ��}�BH���   h�  V�у�P������A  j�� ����4  j ������  ���E�    ��� ���}����  �
��$    �I ��}���   �P����=�  ��  hF  h�  W���Я�����l  j ���E�   �X� ������  h�  W�E�P���Ͱ����}�Q�B<�M��E�7�Ѕ���   V�� ����  �M��L� ������   ����}���   �B����=)  ��   ��}���   �Bx���Ћ�}�Q�Rx�M�Q���҅�uk����� ��p���Q������R3�V�ȉE��� ��tE�������F;�p������4��������I��@;�p���~獅p���P������Q�M�V��� ��u���}���   �P(���ҋ����/������$���j ������0�X  ��}�Q�J�E�P�E�0�ы}����}���   �P(���ҋ��E���<�����$����8 ��   ��}�Q�J�E�P�ы�}�B�Pj j��M�h��Q�҃���}���   ��������R|�E�P�E�8�ҡ�}�H�A�U�R�E�0�Ћ��}�QT3�WP�B�Ѓ�;���  ������Q����� ���}�U��U��M��]�Q�B�PHh�  �������E�9�ҋ�$������������E�0���  �}� ��   ��4��� �E�    ��   3�9s~U��S��}��� ���   �ȋBx�Ћ�$����U������}���   �Bx�Ћ�}�Q�ȋBxW�Ѕ�t1F;s|��s��$����U�<���|jjjV����  ��t�C�<��E�@;�4����E��f�����}�QH�uЋ�p  j h�  V�Ћ�}�QHj �E���p  h�  V�Ћ�}�QH���������   h�  V�Ћ�}�QH�����   h�  V�}��Ћ��� �����(�u�;�t(}+�PV�������  �jj��+�QP�������  3���~5���������d$ ��]�3�;Q��������@����;Ɖ\���]�|ۋ}荅t���P�����������������;�t ��t���}+�PW�  �jj+�WP�  ��}�QH�MЋR8��T���P�ҋ�   �����������P������Q�����R�)�����݅h���3ۃ}�݅`���݅X���݅P���݅H���݅@����  �}�U�����B(����G��    ݅(�����x����H؍t��܅������H������H����]�݅0����H�܅������H������H����]�݅8����H�܅ ������H������H����E���E��Y�Y��x���݅(����L1�H�܅������H���������]�݅0����H�܅������H���������]�݅8����H�܅ ������H���������E���E��Y�Y݅(����H܅������H�����H����x����L��]�݅0����H܅������H�����H���]�݅8����H܅ ������H�����H���E���E��Y�Y��x���݅(����L �H ȃ�`��܅������H������H����]�݅0����H�܅������H������H���ݝ����݅8����H�܅ ������H������H����E��]�݅�������]��E���Y�E��Y�	���;]���   �M��[�D��U�����+�+�݅(�����x����H��ȃ���܅������H������H����]�݅0����H�܅������H������H���ݝ����݅8����H�܅ ������H������H����E��]�݅�������]��E���Y�E��Y�k���������݋���������������;�t&}+�QP�������%  �jj+�PQ�������  �]�3�3Ʌ��y   ���������������<�������u.�r�4��2�������t��r��������t��r��������t���2�4��r��������t��r��������t��������A��;�|���}�B�M���   j j�҅��Y  ��}�HH�uЋ��   j h'  V�ҋ������C  �����������;�t,}+�QP�������  �jj+�PQ�������  �����������;�t&}+�QP��������	  �jj+�PQ��������  ���=� ��ݕ ���3�ݕ���3�ݕ����E�ݕ8���ݕ0���ݕ(���ݕP���ݕH���ݕ@���ݕh���ݕ`���ݝX������e  �d$ ��}�HD�E̋I,�����RWP�ы������v�Ƀ�Ƀ<��:  ��������X������\����T��`����T��d����T��h����T��l����T��������D��@������D����P��H����H��L����P��P����H��T����P�������N�I��(������,����P��0����P��4����P��8����P��<����P�������V�R�Ë�����������X������X������X�� ����X��$����X�������4��������F�D��������]�������������   �������
��@������D����P��H����P��L����P��P����P��T����P�������D��(������,����P��0����H��4����P��8����H��<����P�������N�I������������P������P������P�� ����P��$����P�������4��������V�T���������������4�G;�������M�E�}������SQ�MЍ�t���RPQW������������V��}�P���   j j���Ѕ�t	������N��t����E�"�����ދ�3���}���   �M䋐�   �E���9E��y����M���X 9}�t9{~�UVR��������}�H�A�� ���R�E�!�ЍM�Q�E��sX �U�R�}��E��cX ����  j h���������Y���3�Vhl��M��E�3�E�����}���   �MЋBx�E�4��P�M�Q��t���R�  ������QP��\����5R�]��  P�E�6蚝 ��}�H�A��\���R�]��Ћ�}�Q�J��t���P�E�4�ы�}�B�P�M�Q�E�3�ҡ�}�H�A������R�E�0�Ѓ�,��t����E�"躰����}�Q�J�� ���P�E�!�эU�R�E��TW �u�E�P�E��DW ���M�u��E��R  ������}�B�P�M�Q�ҡ�}�H�A3�Wj��U�h8�R�Ћ�}�Q�J�E�P�E�:�ы�}�B�PWj��M�h,�Q�҃�(��}���   �Bx���E�;��P�M�Q��t���R�  �M�QP��\����<R�]��  P�E�=�6� ��}�H�A��\���R�]��Ћ�}�Q�J��t���P�E�;�ы�}�B�P�M�Q�E�:�ҡ�}�H�A�U�R�E�0�Ѓ�,��t����E�"�Y�����}�Q�J�� ���P�E�!�эU�R�E���U �E�P�}��E���U ��}�}����   ���   �E�P�E��у�������}�H�A������R�Ћ�}�Q�JWj�������h�P�э�����R�E�>�+� ��}�H�A������R�E��Ѓ�������Q�$� ��}���   ���   �M�Q�E��҃��������}��E��CP ��8����E� �4P �������E������"P �   �M�d�    Y_^[��]� ��������̡�}V�񋈈   ���   V�҃��    ^���������������V��V�T ���    ^�������������VW��3�9>t	V�m ���>�~�~�~�~_^�������������U��Q3�9A~V�u�2@��;A|�^]� ���������������U��EV���
�   ^]� �MW��|/�~;�}(�> t#�~ u%��}�H��0  h��h�  �҃�_3�^]� ��;�|���;���_�   ^]� S�;�|�ߋ�+���;ȉ]��   ^��~�F�I���QP�[��P�� ���N��~;ύI�ЉV�'  ������V+ӍR���R��)F+ȍ@��N�N�Q�+�Q贯 �F��}�Q���  �@�h���h�  �PQ�҃������   �N)^�I[��_�V�   ^]� �V��+Ë^�D�����W�@��;ʋ]�E}-�F+�+�����R��R��R�I��R�� �E��;F}L��}�Q���  �@�h���h�  �PQ�҃����u	[_3�^]� �N�I�ȋE�F�V)^[_�   ^]� ��U��EV���
�   ^]� W�}��|/�N;�}(�> t#�~ u%��}�H��0  h��h�  �҃�_3�^]� ��;�|���;���_�   ^]� S�;�|�ً�+���;��]��   ^��~�F��    QP��R�	� ���N��~;ύ��V��   ������V+���R��)F+ȉN�N�Q�+�Q�ƭ �F��}�Q���  h���h�  �PQ�҃������   �N)^[��_�V�   ^]� �V��+ÍD���~��C�^�A�;�}!�U�F+�+���Q׍�Q��R�@� ��;^}C��}�H���  h��h�  ��    RP�у����u	[_3�^]� �V���F�^�])^[_�   ^]� ���U���}�P�B<V���Ћ�}�Q�M�RLj�j�QP���ҋ�^]� �������������U���VW�}���}
_3�^��]� S�]����  �F;ǋ��ύ�N�U��u(��}�H��0  h��h@  �҃�[_3�^��]� ��;���  )^�F�Y  @���j j�и   +�����؋F�ʙÉ]����SP�E��c� �ȉU��;�u��E�;�u�;�|�;M�r��]�Ù9U�E�|�;��{����F�U��NF�@����N��h����u��}�Q���  hV  P�у����}�RhW  PQ��  �у��ȉ�������F�@�F�щN��~N+Ǎ@���P��+E�Í@��P��@��P�� +]��F����Q�[��QP��� ���}  �@�ҋ�+E��R�@���[R��Q�Ҫ ���V  ��~�N����R�@�Q��Q說 ���F�@��ЉN�   �F�D����@����؋F�ʙ;ʉM���   ;���   j jQS�ͭ �ȉU��;������E�;�� ���;E������;�������E�9U�E������;�������h����u%��}�Q���  �[���h{  P�у��$��}�J�[��h|  �RP��  �Ѓ��ȉ���s����F�@�щF�^�F;�}*�N+Ǎ@���R����E�R�@��P�z� ���]�} tG�N;�}"��+��@���R�I�N��j R�H� ���V�[���P���j P�*� ���} tO�N��;�}!�F�I�Ћ�+х�t�P�P�����u�V��ʅ�~�˅�t�P�P�����u��؋E�F[_�   ^��]� ��������������U���VW�}���}
_3�^��]� S�]���  �F;ǋ��ύ�N�U���u(��}�H��0  h��h@  �҃�[_3�^��]� ��;��h  )^�F�.  @���j j�и   +�������F�ʙ��߉}���WS�t� �ȉU�;�u��E�;�u�;�|�;�r��]�Ù9U�|�;�r��M�F�V��Fы���Vh����u��}�Q���  hV  P�у����}�RhW  PQ��  �у�����!����V�}�N���F��~>+�ɋ�+U��QӍ��Q��P�D� �F+]��    Q��RP�,� ���V  �ɋ�+U�Q��Q��R�� ���7  ��~�V��    Q�R��R�� ���F����V�	  �F�D����@����؋F���;���   ;���   j jWS�� �ȉU�;��A����E�;��6���;��.���;��$����E�9U�����;������h����u#��}�Q���  ��    h{  P�у��"��}�Jh|  ��    RP��  �Ѓ����������N���V�^�F9E}"�M�V+���P��P�Eȍ�Q�ԥ ���}�} t=�F;�}�N��+���R��j R誤 ���E�V��    Q��j P莤 ���M��N[_�   ^��]� �������U��j�h9�d�    PQV�Pg3�P�E�d�    �E�    ��}�H�u�QV�E�    �ҡ�}�H�U�AVR�Ѓ���}�Q�B<���E�    �E�   �Ћ�}�Q�M�RLj�j�QP���ҋƋM�d�    Y^��]����������������U��Q�E;�u	�   ]� }+�RP�����]� jj+�PR�����]� ����������U��V��W�~��}_3�^]� jjjW������t�F�M��_�   ^]� �������h�隨 �����U��V���h�脨 �Et	V�cc ����^]� ���������U��M�UV�uW��r�;u��������s��tE��9+�u1��v6�B�y+�u ��v%�B�y+�u��v�B�I+���_��^]�_3�^]�����������U��QV��j �M��;� �F���s@�F�M��O� ^��]�������U��QVW��j �M��
� �G��v	���sH�G�w����֍M�#��� _��^��]�����t�����������U��QW�9��t=j �M�跑 �G��v	���sH�GV�w����֍M�#�軑 ��t
��j����^_��]���̰�������������̸   �����������U��Q�A$V�0W�}j �M�E�    �7�;� �F���s@�F�M�O� ��_^��]� �U��j�hy�d�    PQVW�Pg3�P�E�d�    ���E�    �u���E�    �q�  ��}�H@�Q$VW�E�    �E�   �҃��ƋM�d�    Y_^��]� �����������̡�}�P�B��Q��Y��������������U��MV3���� ��t��}���   ���ȋB(�Ѕ�u��^]� ��������������U��j�h��d�    P��SVW�Pg3�P�E�d�    ���E�    調 �O ���EP�|j P���$� �M�Q���������}�B�P4jh�  �M��E��ҡ�}�P�B4jh�  �M��Ћ�}�E�Q�R8Ph�  �M��ҡ�}�P�B4jh�  �M��Ћ�}�Q@�J(j�E�PV�ы]����3��� ��t&���$    �d$ ��}���   ���ȋB(�Ѕ�u�WV���� ��}���   �Bj j���ЍM��E� ���  ��}�Q�J�EP�E������у��M�d�    Y_^[��]� �����������U��j�hۿd�    P��4SVW�Pg3�P�E�d�    ��u��}�HT�U�Aj R�Ѓ��E��u�M�d�    Y_^[��]� �M�Q���� ���   +��   �]�ƨ   ���Q����������E�    ;�r�h� �N��}�R��i��   �D9 P�BHh�  �M��ЋN+N���Q���������;�r�"� �V��:�    t[S����U  ��}�Q��P�B8h�  �M��ЋM���Q�M���< ��}�B�P<�M�Qh�  �M��E��ҍM��E� �S= �M�E�P�W� �M��E������X�  �   �M�d�    Y_^[��]� ���������������U��j�h.�d�    P��TSVW�Pg3�P�E�d�    ���}��}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�у����   +��   �]�Ǩ   ���Q����������E�    ;�r�� ��}�Q�Rx��i��   G�M�Q���   �ҋ��}�H�A�ލU��R���E������Ѓ�����  ��}�QT�u�Bj	V��3Ƀ��E;�u3��M�d�    Y_^[��]� �MЉM�h�  �M��E�   �� j �M�QP���E�螲 �M��E��� ��}���   �P8�M�Q�҃���uX�E�   �E�   h�  �M��E�跫 j �M�QP���E��e� �M��E�蹝 ��}���   ��M�Q�E��҃��u�E�P��� � S���E��dS  ��}�Q��PP�BHh�  �M���S���BS  ���    t]S���1S  ��}�Q�   P�B8h�  �M��ЋM���Q�M��V: ��}�B�P<�M�Qh�  �M��E��ҍM��E��: �E�P��豿 �M��E���  ��}���   �
�E�P�E������у��   �M�d�    Y_^[��]� ��������������U��j�h��d�    P��TSVW�Pg3�P�E�d�    ���}��}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�у����   +��   �]�Ǩ   ���Q����������E�    ;�r�%� ��}�Q�Rx��i��   G�M�Q���   �ҋ��}�H�A�ލU��R���E������Ѓ�����  ��}�QT�u�BjV��3Ƀ��E;�u3��M�d�    Y_^[��]� �MЉM�h�  �M��E�   �P� j �M�QP���E��ޯ �M��E��R� ��}���   �P8�M�Q�҃���uX�E�   �E�   h�  �M��E���� j �M�QP���E�襯 �M��E���� ��}���   ��M�Q�E��҃��u�E�P���`� S���E��P  ���    t]S���P  ��}�Q�   P�B8h�  �M��ЋM���Q�M��7 ��}�B�P<�M�Qh�  �M��E��ҍM��E��8 �E�P���� �M��E���  ��}���   �
�E�P�E������у��   �M�d�    Y_^[��]� U��j�h��d�    P��TSVW�Pg3�P�E�d�    ���}��}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�у����   +��   �]�Ǩ   ���Q����������E�    ;�r蕠 ��}�Q�Rx��i��   G�M�Q���   �ҋ��}�H�A�ލU��R���E������Ѓ����   ��}�QT�u�BjV��3Ƀ��E;�u3��M�d�    Y_^[��]� �MЉM�h�  �M��E�   ��� j �M�QP���E��N� �M��E�� ��}���   �P8�M�Q�҃���uX�E�   �E�   h�  �M��E��g� j �M�QP���E��� �M��E��i� ��}���   ��M�Q�E��҃��M�E�P�Һ S���N  ـ�   �5���E�   �]�E�]�h  �M��E��� j �M�QP���E�蛬 �M��E��� ��}���   ��M�Q�E��҃�S���M  ���    t]S���M  ��}�Q�   P�B8h�  �M��ЋM���Q�M���4 ��}�B�P<�M�Qh�  �M��E��ҍM��E��5 �M�E�P�� �M��E���  ��}���   �
�E�P�E������у��   �M�d�    Y_^[��]� �������U��j�h7�d�    P��TSVW�Pg3�P�E�d�    ���}��}�H�A�U�R�Ћ�}�Q�Jj j��E�h��P�у����   +��   �]�Ǩ   ���Q����������E�    ;�r蕝 ��}�Q�Rx��i��   G�M�Q���   �ҋ��}�H�A�ލU��R���E������Ѓ�����  ��}�QT�u�BjV��3Ƀ��E;�u3��M�d�    Y_^[��]� �MЉM�h�  �M��E�   ��� j �M�QP���E��N� �M��E�� ��}���   �P8�M�Q�҃���uX�E�   �E�   h�  �M��E��g� j �M�QP���E��� �M��E��i� ��}���   ��M�Q�E��҃��u�E�P���з S���E��K  ���    t]S���K  ��}�Q�   P�B8h�  �M��ЋM���Q�M��(2 ��}�B�P<�M�Qh�  �M��E��ҍM��E��~2 �E�P��胷 �M��E���  ��}���   �
�E�P�E������у��   �M�d�    Y_^[��]� U��j�h��d�    P��  �Pg3ŉE�SVWP�E�d�    ���n ��ݕ������P���ݕ�����������@�Pݝ����������Q������ݕ����R�荅(���ݕ����3�ݝ����P��������d���ݕ���ݕ����ݕ����ݕ(���ݕ0���ݝ8����4}����}�Q�J��0���P�ы�}�B�PVj���0���h��Q�ҍ�0���P�u��| ��}�Q�J��0���P�E������ы��   +��   �����������������X�����	  ��`������   +��   ���������������9�X���r�� ���   �`����{ �   ��x������   ��}�B�P��0���Q�ҡ�}�H�Ij j���x���R��0���P�у���P�����0���R�E�   �[ ��T�����}�H�A��0���R�E������Ѓ���T��� t��T���Q�K� ���U܋E�RP�� ������h������'	  ���   +��   ���������������9�X���r�#� ��}�B���   �P�`���������Q�ҡ�}�H�Aj j�������WR�Ѓ���}���   �R|������P���E�   �ҡ�}�H�A������R�E������Ћ�}�QH���   j h�  V�Ћ�}�QHj ��p������   h�  V�Ѓ��}� ǅt���    ~i3ɍ�    �U�t��d���+���\����t+���l����t�+׉��l���+��p�P��\����P��t���B�� ��;U܉�t���|���h���3�9}���   ��d���݅4���݅L�����p���݅D����R݅<�����ҋ��   ݅�����G��܅�������@܍$��������H��݅����܅�����@܍,��������H��݅����܅����@�������H�����Y��Y��Y�;}�|��������؃; �M  �}� �C  ��E�ݕd���Pݕ\���ݕT���ݕ|���ݕt���ݕl���ݕ����ݕ����ݕ����ݕ����ݕ����ݝ������ ��3҃���l���;���  9U܉�\�����   ��t�������t����M�t
���   �4v�4�V�t
�4v�4�V�t
�L
�4v�I�4���VR��t����x����   ��T���󥋍l���� � ��}�QD��\����R0��T���QVP�҃�t��� F��;u܉�\����i�����l�����h���j W��賷 ��}���   �Bj j����j h�  ���?� ����   ��}�Q�J������P�ы�}�B�Pj j�������hp�Q�҃���}���   �Bx���E�   ��P������Q������R�����P�E��v ��}�H�A������R�E��Ћ�}�Q�J������P�E������у��{ ��  ��}�B�P��@���Q�ҡ�}�H�Aj j���@���h��R�Ѓ����   +��   ���Q��������ʃ����   �E�   ���Qul+��   ��@���R���������u藔 ���   ��}�B����p����H����l���W�ы�}�B��p����PWQ�҃�V���������  +��   �����������  ��@���Q���   +��   ���Q���������u�� ���   ��}�B����p����H����l���W�ы�}�B��p����PWQ�҃�V���G������   +��   ���Q���������   �;��F  ǅt����   h)  �I� ��}�Q������l������&  �J������P�ы�}�B�Pj j�������hd�Q�ҍ�����WP�E���w��P������Q������R�E�������}�Q�R��@���QP�E��ҡ�}�H�A������R�E��Ћ�}�Q�J������P�E��ы�}�B�P������Q�E��ҡ�}���   �R|��<��@���P���ҋ�蓥 3�9u܉�p���~�E�9<�u��p���V�� F;u�|拍h���3��o� ��t$�	��$    ����}���   ���ȋB(�Ѕ�u狍h���V��l���V�Գ ��}���   �Bj j���Ѝ�@���Q���   +��   ���Q���������;�r�ב ��}�Q���   �t������ĉ�p�����p���P�B�Ћ�}��p����Q�JPV�ы�h�����R���������   +��   ��t����   ���Q��������G�;��������h�����}�Q�J��@���P�E������у���P���j j j V���O ��}���   �Pj j����3������������������$����� ��������Ph�   �E�	   �����������ys ���E���������   �M��d��������資 ���   +��   ��X�����`���x��������������F�X���;������   �M�d�    Y_^[�M�3�藃 ��]ËJ��@���P�E������у�3��ʍ�����2� 3����������������U��j�h��d�    P��SVW�Pg3�P�E�d�    �񋎸   +��   ���Q��������3���'  �]����   +��   ���Q���������;�r菏 ���   E��N P��P ����ughG  覡 ��������   ���   +��   ���Q���������;�r�:� ��}���   ���   E��R|P���ҋN j j W�yM WS��� ���WS�������~ W��Su�������1���WS������jj���]� ��}���   �Bj j���Ћ��   +��   �E��   ���Q��������C�;�������   �M�d�    Y_^[��]Ë�}�B�P�M�Q�ҡ�}�H�Aj j��U�h��R�ЍM�Q�E�    �go ��}�B�P�M�Q�E������҃�3��M�d�    Y_^[��]��������U��j�hB�d�    PQSV�Pg3�P�E�d�    ��u����   P�E�   �SE ���   P�GE �����   ��~  ���   3�;�t	P��D �����   P���   ���   ���   ��D ���N\�E��$ �N@�E���# �N$�]���# ��}�H�Q��V�E������҃��M�d�    Y^[��]�����U��j�h��d�    P��SVW�Pg3�P�E�d�    ��u��}�Q�FP�B�Ѓ��N$�E�    �" �N@�E��s" �N\�E��g" ���   ���E��6�  ���   ���E��%�  3��Fx�F|���   ǆ�   �����G�E��E�9Gv�p� ��M��O�M�;Ov�[� �M��U�R�U�RQP�E�P���*g  �{9{v�4� ��M��K�M�;Kv�� �M�U��WRQP�E�P����t  �ƋM�d�    Y_^[��]��������������U��j�h>�d�    P��L  �Pg3ŉE�SVWP�E�d�    ��j��������  �������^\P���E�    ��" ��}�Q�Bdj�������E��Ћ�}�Q�����   h��Gh  W�Ћ�}�Q��jW��`���P�Bh�������Ћ�`���j@jQ�������{�  ��u+�������J���������������y( u��j P��y  ����� ��  ��}�H�A��x���R�Ћ�}�Q�Jj j���x���h��P�ы�}�B�P��h���Q�E��ҡ�}�H�Aj j���h���h�R�Ѓ�(��0���Q���E���! P��h���R�� ���P�E��������x���QP��@����R�]������P�E��Wk ��}�H�A��@���R�]��Ћ�}�Q�J�� ���P�E��ы�}�B�P��0���Q�E��ҡ�}�H�A��h���R�E��Ћ�}�Q�J��x���P�E��ы�}�B�P������Q�E� �҃�4�� ����E��������  �� ���Pǅ ���|��Kt ��3��  ��}�Q�J��h���P�ы�}�B�Pj j���h���h��Q�ҡ�}�H�A��x���R�E��Ћ�}�Q�Jj j���x���h��P�у�(��@���R���E��A  P��x���P�� ���Q�E�	�Y�����h���RP��0���P�E�
�A���P�E���i ��}�Q�J��0���P�E�
�ы�}�B�P�� ���Q�E�	�ҡ�}�H�A��@���R�E����E���}�Q�J��x���P�ы�}�B�P��h���Q�E��ҋ������@��������0������?  �8����������������j
�������z  ��Qh�   ������R��������  j������Ph��Z� �����  ���   ���   ��G��������d����"7  �O���   Q�����  ������R������h��P�� ��}�Q�J��x���P�ы�}�B�@j j�������Q��x���R�Ѓ� �K+K���Q����������E�;�r�� �C�������}�JP�A��x���R�Ћ�}�Q�J��x���P�E��ыK+K���Q���������;�r蹆 �K������Ǆ
�       �  j������Ph���#� ����uJ���   +��   ���Q���������;�r�`� ���   �DP������h��Q踒 ���Q  j������Rh��迒 ����uJ���   +��   ���Q���������;�r��� ���   �TR������h��P�T� ����  j������Qh���[� ����uJ���   +��   ���Q���������;�r蘅 ���   �TR������h��P�� ���  j������Qh|���� ����uC���   W���4  ��0PW���	4  ��(PW����3  �� P������hl�R蓑 ���,  j������Phh�蚑 ����uC���   W���3  ��HPW���3  ��@PW���3  ��8P������hX�Q�6� ����  j������RhT��=� ����uC���   W���[3  ��`PW���O3  ��XPW���C3  ��PP������hD�P�ِ ���r  j������Qh@���� ����uC���   W����2  ��xPW����2  ��pPW����2  ��hP������h0�R�|� ���  j������Ph(�胐 ����uZ������Q������h�R�B� ��j ������P������@Q�������Q���   W���E��g2  �ȃ��h��������yj������Ph��� ������   ������Q������h�R�ʏ ��j ������P�� �����P���� ���Q���   W���E���1  �ȁ��   �g���� �����}�B�PQ�E��҃�W���1  ǀ�      �������@������������������l  ��u+�������I���������������y( u��j P�q  j��d�����  ��T����^@R���E��� ��}�P�Bdj��T����E��Ћ�}�Q�����   h��Ghd  W�Ћ�}�Q��jW��`���P�Bh��T����Ћ�`���j@jQ��l����b�  ��u+��d����J��l�����d������y( u��j P��p  ������ ��}�H�A��h���R��  �Ћ�}�Q�Jj j���h���h��P�ы�}�B�P��x���Q�E��ҡ�}�H�Aj j���x���h�R�Ѓ�(��@���Q���E�� P��x���R�� ���P�E��������h���QP��0����R�]�����P�E��>b ��}�H�A��0���R�]��Ћ�}�Q�J�� ���P�E��ы�}�B�P��@���Q�E��ҡ�}�H��x����E�R�A�Ћ�}�Q�J��h���P�E��ы�}�B�P��T���Q�E��҃�4�������E���}  �������|�P�������4k ��}�Q�J������P�E� �у��� ����E������}  �� ���R�� �����j ��3���  �Ћ�}�Q�Jj j���h���h��P�ы�}�B�P��x���Q�E��ҡ�}�H�Aj j���x���h��R�Ѓ�(��@���Q���E��� P��x���R�� ���P�E�������h���QP��0����R�]������P�E��` ��}�H�A��0���R�]��Ћ�}�Q�J�� ���P�E��ы�}�B�P��@���Q�E��ҡ�}�H��x����E�R�A�Ћ�}�Q�J��h���P�E��ы�d����B3���0��l�����������  j
��d�����p  ��Ph�   ������Q��d����݈  ���   +��   ���Q��������3����   ��d�����}�Q�J��x���P�ы�}�B�@j j�������Q��x���R�Ѓ����   +��   ���Q����������E�;�r�~ ��}�B���   �d����@x��x���R�Ћ�}�Q�J���ߍ�x����PG�E��у���u2���   +��   ��d����   ���Q��������C�;��&����������������j������Qh���� �����,  ���   +��   ���Q���������;�r�M} ���   i��   ���   R������h��P蜉 ��d����I��j
��d����'o  ��Rh�   ������P��d����,�  ��}�Q�J��h���P�ы�}�B�@j j�������Q��h���R�Ѓ����   +��   ���Q����������E�9�����r�| ���   ��}�H�A���   ��h���WR�Ћ�}�Q�J��h���P�E��ы�������   j	������Rh���ʈ ������   ��d����Hj
��d����+n  ��Qh�   ������R��d����0�  ��}�H�A��P���R�Ћ�}�Q�Rj j�������P��P���Q�҃����   +��   ���Q����������E�;�r�{ ���   ��i��   ���   ��}�Q�JP��P���P�ы�}�B�P��P���Q�E��҃���d����@��l����k���3���l���9�����t ���V  ��u3�������Q�m� ����t3���t�����|�����x�����������������������������������}������������ƅ���� ƅ���� ��������������x�����������������t���������������������������������;�u)��d����H��l�����d�����9y(u��WP�0i  ��`���V�� ������Y  ��}�Q�J�����P�ы�}�B�PWj������h��Q�ҡ�}�H�A�� ���R�E��Ћ�}�Q�JWj��� ���h�P�ы�}�B�P��P���Q�E��ҡ�}�H�AWj���P���VR�Ѝ�P���Q�� ���R������P�E� ������H�����QP�������!R�]������P�E�"�|Z ��}�H�A������R�]��Ћ�}�E� �Q�J������P�ы�}�B�P��P���Q�E��ҡ�}�H�A�� ���R�E��Ћ�}�Q�J�����P�E��у�$��}�B�P��T���Q�E��҃��������E��$v  �������|�P�������oc ��}�Q�J������P�E� �у��� ����E�������u  �� ���R�� ����/c ���   �M�d�    Y_^[�M�3��k ��]����������V���8����������   ^�����������U��j�h��d�    P��$SVW�Pg3�P�E�d�    3��u�M�u��X�  �E�]jV�M�Q�ˉu��E�   �E���7  �������   �U�U��    ��+�PV�M�Q���Z  �MP�E�   �ϋ  �}��E� r�U�R�. ��j�wV�EP���x7  �����u�PV�M�Q���tZ  �uP���E�   肋  �}�r�U�R�c. ���ƋM�d�    Y_^[��]� �E�M�d�    Y_^[��]� ���U��j�hJ�d�    P��  �Pg3ŉE�SVWP�E�d�    �u�ٿ   W��������~  j@WV�������E�    ��v  ��u+�������H���������������y( u��j P�Ge  ��8��� ��  ��}�Q�J������P�ы�}�B�Pj j�������h��Q�ҡ�}�H�A��p���R�E��Ћ�}�Q�Jj j���p���h�P�ы�}�B�P������Q�E��ҡ�}�H�Aj j�������VR�Ѝ�����Q��p���R������P�E��!�����H������QP������R�E�����P�E��V ��}�H�A������R�E��Ћ�}�Q�E��J������P�ы�}�B�P������Q�E��ҡ�}�H�A��p���R�E��Ћ�}�Q�J������P�E� �у�$��<����E������\r  ��<���Rǅ<���|��_ ��3��k  ��}�H�A������R�Ћ�}�Q�Jj j�������hT�P�э�����R�E��V ��}�H�A������R�E� �Ћ������A������������  j
�������Xf  ��Rjc������P�������`~  j������QhD�誀 ����uK{|���   +��   ���   ���������������;�r��s ���   ����+�|�h�D�h�!  j������PhP��E� ����uN��   ���   +��   ���   ���������������;�r�ts ���   ����+�|�l�D�l�  j������Qh���� �����  ��   ���   jx������@j R�������j ��l���   ������󥋍�������   Q���q  ���   +��   ���   ���������������;�r��r ���   ����+�3��|�d���   +��   ���   ���������������;�r�r ���   ����+Ή|�h���   +��   ���   ���������������;�r�Er ���   ����+Ή|�l�   �  j������PhL��~ �����k  {x�������������   �������������P���@��u�+�P������Q�������H  WW������R��P����E��{  �������E�	r������P��( ��������������ǅ����    ƅ���� ���  ������Q�� ���     �p�@    �������@ �� ��P����̉�����R�E��=�  ������P�E�
��  ������+�������$I�����������t
���H����   t#��t~3���   R���   �e  ��d���0����   P���   �I  ��d8�������Yt  ��P����E� �@  �������A�������=����������8Z  ��u+�������J���������������y( u��j P�9_  �{|3ɋǺ   �������Q�~& �����������E�����   h�$ WjV�>����   ��}�B�P������Q�ҡ�}�H�Aj j�������h4�R�Ѝ�����Q�E���P ��}�B�P������Q�E�
�҃��������Ks  �������E� ��6  �������|�P�������WZ ����<����E�������l  ��<���Q��<����0Z ��3���  3����   3ɋǺ   �����E� ���   ���Q�j% �����������E���th�$ WjV�=���3����   ���   +��   ��������������3���E� �C  3����   +��   ���������������;�r�n ���   ǋ@d3�@�    �������Q��$ ���   +��   ���������������������;�r�Nn ���   �������Tp���   +��   ���������������;�r�n ���   ǋ@d3�@�   �������Q�=$ ���   +��   ���������������������;�r��m ���   �������T9t���   +��   ��������������F�x;��������<����E�������j  ��<���Qǅ<���|��;X ���   �M�d�    Y_^[�M�3��` ��]� ���U��j�h��d�    P��  �Pg3ŉE�SVWP�E�d�    �]��������������|�  3��������u��l�  j�������E��+u  j@jS�������E��m  ��u)�������H��������������9q(u��VP�z[  9�������  ��}�Q�J������P�ы�}�B�PVj�������h��Q�ҡ�}�H�A�����R�E��Ћ�}�Q�JVj������h�P�ы�}�B�P��t���Q�E��ҡ�}�H�AVj���t���SR�Ѝ�t���Q�����R��@���P�E��X�����H������QP��(����R�]��<���P�E���L ��}�H�A��(���R�]��Ћ�}�E��Q�J��@���P�ы�}�B�P��t���Q�E��ҡ�}�H�A�����R�E��Ћ�}�Q�J������P�E��у�$�������E��h  ������Rǅ����|���U ���������n  �������n  3��s  ��}�H�A�����R�Ћ�}�Q�JVj������h��P�ы�}�B�P��t���Q�E��ҡ�}�H�AVj���t���h��R�Ћ�}�Q�J������P�E�	�ы�}�B�PVj�������SQ�ҍ�����P��t���Q��(���R�E�
躼����H�����QP��@����R�]�螼��P�E��4K ��}�H�A��@���R�]��Ћ�}�E�
�Q�J��(���P�ы�}�B�P������Q�E�	�ҡ�}�H�A��t���R�E��Ћ�}�Q�J�����P�E��ы�}�B�P��l������Q�������������ҡ�}�H�A������R�E��������Ћ�}�Q�JVS������h��P�э�����R�E��<K ��}�H�A��������@R�E��Ћ������A������������  3�ǅ�����������������������$    �d$ j
��������Z  ��Rh�   ������P��������r  j������Qh���!u ������   ������R������h��P��t �������Q��P����,�  ��P����w\R���E�� ��P����E����  ���Q ������P��P������  ��P���Q���E�� ��P����E���  �  j������Rh���st ������  ��}�H�A��t���R�Ѓ��������������E�������;�v�g ��������������������;�v�g ������������QSVR�����P�������m  ������ǅh���   ǅd���    ƅT��� �P���@��u�+�P������Q��P����d=  jj��P���R��l����E��Zp  ��h���r��T���P�5 ��������P3҃� �Ĺ   ��H�P��h�����d�����T����������P�� ��l����̉�����R�E��y  ��|���P�E��q|  ������������+θ�$I����������ʃ�H��w�Zf �������~4r�v ��� ��}�B�P������Q�ҡ�}�H�Aj j�������VR�Ћ�}�Q�R��t���P������Q�E��ҡ�}�H�A������R�E��Ћ��   +��   ���   ���Q���������� 3��t{���������$    �N+N���Q���������;�r�e ��}�B�N������@x��t���R�Ѕ��  �N+N�������   ���Q��������C�;�r��N+N���Q�������   ���̍\�������  S���@d  �N+N���Q��N+N������ڸ��Q��������K�;�r��d ��}i��   ^�B�P��t���SQ�ҋN+N���Q���������L��������������E���+  ������Rǅ����|��DO ��}�H�A��t���R�E��Ѓ���  �������j������Qh����p ����u@������������x@P���   �������������  P������h��R�cp ���z  j������PhD��jp ����u8���   ��������HQ�PRP������h��P�p ���������(  j������QhP��p ����ud���   ��HQP������h��R��o ���   ÍHQ�PRP������hx�P�o �苏�   �d�D��$����������  j������RhL��o ������  ���������t������P���   �e  �Ht����������������j  ������P��P����E  jj��P���Q��l����E���k  ��P�����2  ������R�� �ĉ0�@   �p�������@ �� ��l����̉�����P�E��Zu  ��p���Q�E��*x  ��H�������<j  ������+�������$I�����������T����������x  ���o  �  ��8����������m�  �� ����E��^�  �   �E�9������  j/S�������  P��T���Q������P�������E��o  ��T����E��-e  j �������  �xr�@���P�n ����������NR��8����������Ne  h��j�������<  P�2  ����t=j�������"  �xr�@���P�[n H��������������P�� �����d  ���   �v�D��ʋ���������\$�@�\$� �B�$��C;�����������������p���R����l����$P�҃�l��� ������ǅ����    �f  ��H���ǅ����    ���    3۹   +˃�u3ɋ�����+�D���ы������4�����������;�r�` ���   +��   ��D����4����������������9�����r��_ ���������   �ˋ������Dp�����H�����+�D�������vz��0���+�,����������0��;�r�_ ���   +��   ��,����4����������������9�����r�^_ ���������   �ˋ������Dp��L���H���C�������������������������A������;�l��������������R�Vy  ��,���3���;�t	P�1 ���� ���P��,�����0�����4���� ��D�����;�t	P�� ����8���Q��D�����H�����L����� ����  ǅ����   ���  ������������I ������j/R�������\  P��T���P���=���P�������E��=l  ��T����E���a  j �������!  �xr�@���P�Zk ��������Q���   �X��u  �Pph��j�������\2���  P�F/  ����t@j��������  �xr�@���P��j �X���������P���   �  �Hp�\1������@��������;�����������������   j �������Y  �xr�@���P�j ��������������H���   R�ˉ��������  �@p������h���L0j��������  P�i.  ����tFj��������  �xr�@���P�j ��������HR�ˉ������9  �@p�������L0�������������E���#  ������Rǅ����|��SG ��������3��������@�����������������9�����t ���7  ��u3�������Q�g ����t3���������������������������������������������������}������������ƅ���� ƅ���� ������������������������������������������������������������������;�u)�������H��������������9q(u��VP�PJ  ��}�Q�J��l���P�E��у��������E��X  ������Rǅ����|��F ��������;�t*��p���Q������������RQP�H  ������R�; ��������P������������������� ��������;�t*��p���Q������������RQP�RH  ������R�� ��������P�������������������� ���   �M�d�    Y_^[�M�3��M ��]� ���������������U��j�h�d�    P��<  �Pg3ŉE�SVWP�E�d�    �E�}��F ��}�Q���   j j	���Љ��}�Q���   j j���ЉF��}�Q���   j j���ЉF��}�Q���   j j
���ЉF��}�Q�J������P�у�������Rj������P���E�    �J'����}�R�NQP�B�E��Ћ�}�Q�J������P�E� �ы�}�B�P������Q�E������ҡ�}�H�A������R�Ѓ�������Qj������R���E�   ��&��P�������E����  �������^$P���E��T�  �������E��U�  ��}�Q�J������P�E��ы�}�B�P������Q�E������҃�h���������M�  ������P���E�   ��  �������E��������  ��}�Q�J������P�у�������Rj������P���E�   ��%��P�������E�� �  �������~@Q���E��{�  �E��������|�  ��}�B�P������Q�E��ҡ�}�H�A������R�E������Ѓ�h���������u�  ������Q���E�	   �0�  ����������}���  j��������_  ������R���E�
   ��  ��}�Q�Rhj h�   ������Q���E��ҡ�}�H�A������R�E�
�Ѓ�j@j������Q�������ZW  ��u+�������J���������������y( u��j P�E  ����� ��}�H�A�V  ������R�Ћ�}�Q�Jj W������h��P�ы�}�B�P������Q�E��ҡ�}�H�Aj W������h�R�Ѓ�(������Q���E���  P������R������P�E�軨��������QP��d����R�]�袨��P�E��87 ��}�H�A��d���R�]��Ћ�}�Q�J������P�E��ы�}�B�P������Q�E��ҡ�}�H�E��A������R�Ћ�}�Q�J������P�E�
�у�0������}���R  �����Rǅ���|��I@ ��3��  ������R�Ћ�}�Q�Jj W������h��P�ы�}�B�P������Q�E��ҡ�}�H�Aj W������h��R�Ѓ�(��d���Q���E��M�  P������R������P�E��e���������QP�������R�]��L���P�E���5 ��}�H�A������R�]��Ћ�}�Q�J������P�E��ы�}�B�P��d���Q�E��ҡ�}�H�E��A������R�Ћ�}�Q�J������P�E�
�ы������J��0j
�������>F  ��Ph�   ������Q�������C^  �������=  ��u+�������J���������������y( u��j P�B  ������P�_ ��;��`  ��}�Q�J������P�ы�}�B�Pj W������h��Q�ҡ�}�H�A��t���R�E��Ћ�}�Q�Jj W��t���h�P�ы�}�B�P������Q�E��ҡ�}�H�Ij W������R������P�э�����R��t���P��T���Q�E�膥����H������RP��D����P�]��j���P�E�� 4 ��}�Q�J��D���P�]����E���}�B�P��T���Q�ҡ�}�H�A������R�E��Ћ�}�Q�J��t���P�E��ы�}�B�P������Q�E�
�҃�$�=4 ������P���_���������Q�������~ t-���   +��   ���Q���������t���%�������������g�����3 j h  �4 ��������}��UO  �����Qǅ���|��< ���   �M�d�    Y_^[�M�3���D ��]� ���������Q�|��f< Y��̋A��P�D
�����U��V��N+N��������������W�}�;�r�KQ �V����+�_��^]� �U��V��N+N���Q��������W�}�;�r�Q ��i��   F_^]� �����U��V��N+N��$I����������W�}�;�r��P �V��    +�_��^]� ���������������U��V��蕥���Et	V�� ����^]� ���������������U��j�hb�d�    PQV�Pg3�P�E�d�    ��u��}�H�QV�����V0���   �V(P�V �E�    �VH�V@�V8�V`�VX�VP�Vx�Vp�^h��}�Q�B�Ћ�}�Q���   P�B�E��Ћ�}�Q���   P�B�E��Ћ�}�Q�J���   P�E��у��ƋM�d�    Y^��]��������U��j�hb�d�    PQV�Pg3�P�E�d�    ��u��}�H�A���   R�E�   �Ћ�}�Q�J���   P�E��ы�}�B�P���   Q�E��ҡ�}�H�A���   R�E� �Ћ�}�Q�BV�E������Ѓ��M�d�    Y^��]����������U��V��V�|��9 ���Et	V�� ����^]� �����U��A�U��Q �E��U+ЋA0�]� ��������������̋A �8 t�I0��3�����������������U��A�U��Q$�E��U+ЋA4�]� ���������������V���F@t�F�Q�\ ���V�    �F �     �N0�    �V�    �F$�     �N4�    �f@��F<    ^�������U��Q�A8V�0W�}j �M�E�    �7�k4 �F���s@�F�M�4 ��_^��]� ̍Q�Q �Q�Q$�A�A�Q(�Q0�A�A�Q,�Q4�     �A$�     �Q4�    �A�     �Q �    �A0�     ���������U��j�h��d�    PQSVW�Pg3�P�E�d�    ��u��}�H�QV�ҡ�}�H�}�QVW���G�^���   �GS�^�G�F�O �N �W$�V$�G(�F(�O,�N,�W0�V0�G4�F4�O8�N8�W<�V<�G@�F@�OD�ND�WH�VH�GL�FL�OP�NP�WT�VT�GX�FX�O\�N\�W`�V`�Gd�Fd�Oh�Nh�Wl�Vl�Gp�Fp�Ot�Nt�Wx�Vx�G|�F|��}�Q�B�E�    �Ћ�}�Q�J���   SP�ы�}�B�H���   S�E��ы�}�B�P���   SQ��ه�   ٞ�   ��}�H�Q���   S�E��ҡ�}�H�A���   SR�Ћ�}�Q�B���   S�E��Ћ�}�Q�J���   SP�ы��   ��<���   �ƋM�d�    Y_^[��]� �����U��VW�����u�5K ���t��3ҋE����+��G����;Bw��t�	�3�;As��J w��_^]� ���������U��VW�����u��J ���t��3ҋE�4�    +��G���;Bw��t�	�3�;As�J w��_^]� ���������U��M����w3ɋ���+����R��  ����]Ã��3����xsڍEP�M��E    ��E h�;�M�Q�E�h��:J ���U��M����w3�i��   Q�U�  ����]Ã��3���=�   sߍEP�M��E    �E h�;�M�Q�E�h���I ��������U��M����w3ɍ�    +���R���  ����]Ã��3����sڍEP�M��E    �-E h�;�M�Q�E�h��zI ���U��M����w3ɍ�    R��  ����]Ã��3����s��EP�M��E    ��D h�;�M�Q�E�h�� I ���������U��EVP����D �h���^]� ����U���}VW�}��H�QVW���G�^�G�^�G�F�O �N �W$�V$�G(�F(�O,�N,�W0�V0�G4�F4�O8�N8�W<�V<�G@�F@�OD�ND�WH�VH�GL�FL�OP�NP�WT�VT�GX�FX�O\�N\�W`�V`�Gd�Fd�Oh�Nh�Wl�Vl�Gp�Fp�Ot�Nt�Wx�Vx�G|�F|��}�Q�R���   P���   Q�ҡ�}�H�I���   R���   P��ه�   ٞ�   ��}�B�@���   Q���   R�Ћ�}�Q�R���   P���   Q�ҋ��   ��(���   _��^]� ���U��S�]V�u;�t#W�}V���������   ���   ;�u��_^[]ËE^[]��������U��S�]V�u;�t#W�}���   ���   V���I���;�u��_^[]ËE^[]��������U��E��V��M�Q�F����- ��V�H�N�P�V�@�F����^��]� ���������������U���E��QP�+ ��]� ��������U��S�]V�u;�tW�y�WP�+ �F��;�u�_��^[]� U���E��QP��1 ��]� ��������U��S�]V�u;�tW�y�WP�1 �F��;�u�_��^[]� U��E]� ������U��E�UV�1W��+�W�}WP�FR��_^]� �������������U��S�]VW�}��+�9us��E �E�MVSPQ��B ����_^[]� �����������U��E]� ������U��E�UV�1W��+�W�}W�}WP�F(R��_^]� ���������U��S�]VW�}��+�9us�ME �E�MVSPQ�MB ����_^[]� �����������U��V��F�����~�FP�gE �}�NQ��  ���E�t�t	V�2�  ����^]� ��������V��W�~8�����t��踙��W��  ��_�N^��/ ����̃��� ����������3��������������̃���������������U��U��@R�Uj�R��]� �������̋�� ������������ ������������̋A$�8 t�I4��3�����������������V���P�҃��u�^ËF0��F ��Q��^����������U��E�x��3ɉH�H�H]� ���U��E�x��3ɉH�H�H]�  ���U��A � ��t<�Q;v5�U���t:P�t�A@u"�A0� �A ����t�A ����]� 3�]� ���]� ̋Q V�2��u���^�SW�y0����;�s�_[^��A@u/�A$� ��t&;�w9q<v9A<s�A<��A<+�I ��_[^�_[���^����������������U��SV�q$�W��t9A<s�A<�]����   �A �����   �E��u�A�y<+8�u��'��u��u�A�u��+8����t�5x���u����   �A� �y<+�;���   +Q0�)�Q ����   �Q$�����   �Q4�ЋA R��AR�R������p��te���t_�E�=x���u�A�Y<+�u����u�A�u��+��	����u�u��|�A� �Y<+�;�+Q4�)�I$�
����5x��E_3ɉ0^�H�H�H[]� ��U��E�UVW�y$�4���t9A<s�A<�x�;���   S�]$��tR�Q ���tI��|w�A� �y<+�;�d+Q0�)�Q ��tX�Q$���tO�Q4�ЋA R��AR�R�����4��t-�?��t'��|#�A� �Q<+�;��Q4+��)�I$��x���[�E3�_�0�H�H�H^]�  ��������������U��V�q���Q�F�D���P� |��o+ ���Et	V���  ����^]� ����U��V��W�~8�����t���U���W��  ���N�|+ �Et	V��  ��_��^]� �������������U��V��W��������~8�����t�������W�D�  ���N�!+ �Et	V�-�  ��_��^]� ��U��Q�U�E�M���u	;A��   SVW�y;�st+�;�wn�   +���yr
���M�	����M��E�WQS�= ������t5�U�ERPV�_�������t,�M�+ލ|�WR�^S��< ������u�_^���[��]� �E��x�Mr�	_��^+�[��]� �U��SV�uW��9ws��+ �G+Ƌu;�s���]��;�r�Ãr�����MP�EP�W�Ē������u;�s
_^���[]� 3�;���_^[]� �U��M����w3�Q���  ����]� ���3����s�EP�M��E    �: h�;�M�Q�E�h��e> ��������������V�����t(��u�4> ��xr�H��H�@�9Fr�> �F^����������U��E��u&�yr�I�E�U�]� �E�U���]� �yr�I����UP�EP�Q�4 ��]� ���������U��j�h��d�    P��SVW�Pg3�P�E�d�    �ى]�K����( j�E�    ��  ������t.��& ���$ j �M����$ �G���s@�G�M��$ �3��ˉs8�����ËM�d�    Y_^[��]�U��S�]V�uW���    ��t)��t%�V�F��r����;�w��r� �N�;�v��< �7�_��_^[]� ������������U��E�M�UV�uPQRV�9 ����^]����������������U��E�M�U ��E��   ]� ����U��E�M��   ]� ������������U��E+E�M;�s��]� ����������U���EV���t�t	V�H�  ����^]� ��������������U��S�]V�u��+θ����������������+ȋE�ȉM��;�t#+�W��I �<���x�   �;�u�E_^[]�^��[]����������������U��S�]V�u��+˸����������������+���ɋыM��+�;�t+�W�M��M��x�<�   ���;�u�_^[]����������������U����US�]V�uW�}2��E��M��E��E�PQRWVS����+���Q���������i��   ����_^+�[��]����������U��U�ES�];�tVW��t�   �����x��x;�u�_^[]���������������̋��Q�D(��t�H�% ���������V��F � ��t=�N0�	��~�F0��F � �V �� ^Å�t�N0�9 ~����F ��Q���	��P���҃��u�^ËF �8 t�N0�9 ~��^Ë�P��^������U��QV3�9uW���u�~nS�]���3�����~6�M;ȋ�}��G ��UVQRS�6 �G0)0u�)u�G ރ�0�u����P���҃��tF�C�M�u��} �[_��^��]� _��^��]� ������U��QV3�9uW���u�~mS�]���������~3�M;ȋ�}��VSP�G$�Q�6 �G4)0u�)u�G$ރ�0�u����P�B���Ѓ��tFC�M�u��} �[_��^��]� _��^��]� �������U��j�h�d�    PQVW�Pg3�P�E�d�    �M��A��P�D
����q����E�    ���3����~8�����t���?���W��  ���N�f# �F��H�D1����M�d�    Y_^��]����������������U���V���F@Wt �~$���t�N<;�s�F4� +��N4��E���u
_3�^��]� �V$�:S��t$�N4����;�s�	�v$�[�Q�_�^��]� �F@u=��u3���F4�N�+ߋ���� s�    ���v������+�;�s��u��u[_���^��]� �P�ND�E��������F��M���vSQ�M�QW�y����M�����u"�V�~<�:�F$�8�V4�E���F@u7�GPW�V�F$��+�V<� �V��+�+��V$ǉ��+�U��F4��F@t�V�:�F �     �V0�:��F$��F BR�+��RW��������M��F@t	Q���  ���F4�N@��v$��A��E[_�^��]� �����������̋P��  Y�������U��S�]V��W9^s�%# �F�}+�;�s����v^�N��r�V��V�U��r�V��V+�P�E��P+�Q�R�04 �F+ǃ��~�Fr�N_� ��^[]� �N� _��^[]� ��U��} VW�}��t'�~r!�FS���vWSjP�2 ��S���  ��[�~�F   �D> _^]� ����U��E�MPQ�D7 3҃������]�V��~L t#��Pj��҃��t�FLP�; ����}���^�3�^�U��A � S�]��t,�Q9s%���t�@�;�u�A0� �I �	��@���#�[]� �AL��t$���t�y< u��PQ�8 �����t��[]� ���[]� �V��F ���t�Ћ�V0��;�s�^Ë�PW���ҋ����u_�^Ë�PW���ҋ�_^������������U��V��NLW��tl�U�}��u	��u�G�3�WPRQ�n: ����uG�~L���FH�FA������t�G�F�F�G�~ �~$�F0�F4�~L��}�FD_�F<    ��^]� _3�^]� ��������������U��ES�]V���F<    �F@����   ��<tzWS�ND��������ESPSW�0 ���F@��F<u�N�9�V �:�N0��N@��u7��u�ǋV�:�N$���+ЋF4Ӊ�N �9 u�V�:�F �     �N0�9�N@_^[]� ����������U��V�1W�y��u�3 3��Mi��   �;xw��t�����3�;xs��2 �E�x_�0^]� �����U��j�h0�d�    P��SVW�Pg3�P�E�d�    �e����}�E�������v���"�_������������;�s�����+�;�w�4�NQ���E�    �����E�&�E�M�E�@�e�P�E������E�zË}�u�]��v �r�G��GSP�E�VRP�/ ���r�OQ�:�  ���M�G�  ��w�_��r��� �M�d�    Y_^[��]� �u�~r�VR���  ��j �F   �F    j �F �1 �������U����US�]V�uW�}2��E��M��E��E�PQRWVS�����+���Q���������i��   ���_^[��]��������������U��E�U;�tS�]VW����x�   ���;�u�_^[]�������U��V�uW�};�tS�]S����������   ;�u�[_^]�������U��U��v#�ES�]VW��t�   ����J��x��w�_^[]��U��j�ha�d�    P��SVW�Pg3�P�E�d�    �e��u�}3ۉu�]���$    ;}tU�u�u��E�;�tW���������   �]��u���   �ыu�};�t��$    ���y������   ;�u�3�SS�0 �ƋM�d�    Y_^[��]���V�qP���5���V�|�� ��^�����V��~r�FP���  ��3��F   �F�F^�����������U��VW�y��wP�������V�|��T ���Et	W��  ����_^]� ��������U��yr�AV�uQP���7�����^]� V�u�AQP��� �����^]� ���������U��j�h��d�    PQV�Pg3�P�E�d�    ��u��B����E3ɉM����u�   �u���t���t���E�x�Pr�@���QRP��������ƋM�d�    Y^��]� ����U��U��V�p�d$ �@��u��M+�P�ARPj �G��������^]���������������U��Q�M�U�E� �E�P�EQ�MR�UPQR��������]�����U��Q�M�U�E� �E�P�EQ�MR�UPQR���������]�����U��j�h��d�    P��SVW�Pg3�P�E�d�    �e��u�}3ۉu�]���$    ;�vL�u�u��E�;�t�EP���c���O���   �]��u�ԋu�};�t����������   ;�u�3�SS�g- �M�d�    Y_^[��]���������������V�����~$r�FP�h�  ��3��F$   �F �F��^�c) �������������̃y$r�AÍA���U��j�h�d�    PQSV�Pg3�P�E�d�    ��u�3�S�z �   �F�^�]��^�F8�^4�^$�FT�^P�^@�Fp�^l�^\�EPV�E�� ���ƋM�d�    Y^[��]� ������������U��j�hd�d�    PQSVW�Pg3�P�E�d�    ��u�V�E�   �� ���~pr�F\P�V�  ��3ۿ   �~p�^l�^\�~Tr�F@P�4�  ���~T�^P�^@�~8r�F$P��  ���~8�^4�^$�~r�FP���  ���~�^�Έ^�E������ �M�d�    Y_^[��]���V��~r�FP��  ��3��F   �F�F^�����������U��S�]V�����+F;�w�� ����   W�~����v�� �F;�s9�NQW���L�����vZ�U�FRSP��������~�~r:�F�8 _��^[]� ��uщ~��r�F_�  ��^[]� �F_�  ��^[]� �F�8 _��^[]� �����U��S�]VW�}��9_s� ��E+�;�s���M;�uj��W���'���Sj ������_��^[]� ���v� �M�F;�s�FPW���t����M��vj�yr/�I�-��u�~��r�F_�  ��^[]� �F_�  ��^[]� ���~�^r���ËUW�Q�NQP��& ���~�~r��; _��^[]� ����������U��USVW���tF�~�F��r����;�r1��r���ȋ^�;�v��r� �MQ+�RV�������_^[]� �}���v� �F;�s�VRW���{�����vY�N�^��r.��,��u�~��r�F_�  ��^[]� �F_�  ��^[]� �ËUWRQP�& ���~�~r��; _��^[]� �����U��Q�UV�uW�}�E� �E�P�ER��QPVW������΃���+΍�_^��]� ����U��V3���j��F�F   P�F�EP�������^]� ��������U��j�h��d�    P��D�Pg3ŉE�SVWP�E�d�    �A � 3҉M�;�t'�A �q0� �6�;�s�A0��A ��Q���K  �AL;��=  9Q<uP��( ������&  ���!  �E�   �U�U�P�U��( �������  Pj�M��Y����}�E؃��5  ���u̅�t!�ȃ�s�M�;�w�ȃ�s�M؋U��;�v�r' �}�U�E؍Mԃ��t�ȃ�s�M��;�r�L' �}�U�E؋ڃ���   ����t�ȃ�s�M�;�w�ȃ�s�M��;�v�' �}�U�E؍Mԃ��t��s�E��;�r��& �}ċO<��R�E�P�E�P�E�P�E�P�E��PV�GDP�҅���   ��~_����   �}���   j�U�R�M��>������G���P�E�jP�# �uӃ��M��������   �M؉M̋�������u��%����E�9E���   �U�E؃���   ����t!�ȃ�s�M�;�w�ȃ�s�M؋]��;�v�& �U�E؍Mԃ��t��s�E؋U��;�r��% �E�+�Pj �M������OLQ�& ����������M����������M�d�    Y_^[�M�3��� ��]Íu��b����}�M�Q�M��2������;���+}ȋ����~�UċBL�M��T�NPR�L) ������uӍM�����������U��V�u��W�x�I �@��u�+�PV�p���_^]� ����������U��SVW�}���    ��t�E9Fw;Fv��$ �E�]���G9^w;^v��$ �]����t;�t��$ �O;�t!�F�E �UR�UR�URQPS�������F��_^[]� ��������U��j�h��d�    P��,�Pg3ŉE�SVWP�E�d�    �y< �M���  �yA ��  ��Pj��҃���m  �   3��E� �M�E؉E��E�   ��s�E��@ �E�    �E؋U����    ����   �؉]̅�t!�ȃ�s�M�;�w�ȃ�s�M؋u��;�v�# �U�E؍Mԃ��t�ȃ�s�M؋u��;�r�# �U�E؋}����   ����t$�ȃ�s�M�;�w�ȃ�s�M؋]�ˋ]�;�v�X# �U�E؍Mԃ��t��s�E؋U��;�r�4# �EЋH<��R�E�P�E��SV��DP�҃� t)��t+���M��7  �>  �]؉]������u��i����E��@A �U�E؃���   ����t!�ȃ�s�M�;�w�ȃ�s�M؋}��;�v�" �U�E؍Mԃ��t�ȃ�s�M؋}��;�r�" �U�E؋}�+�tv����   ����t!�ȃ�s�M�;�w�ȃ�s�M؋]��;�v�@" �U�E؍Mԃ��t��s�E؋U��;�r�" �EЋHLQWjV�* ��;�u7�U�E؋MЀyA t4�������Wj�M�����������u������u��h����M������2��
�M��������M�d�    Y_^[�M�3��� ��]������U��V�uW�};�t�����������   ;�u�_^]� ���������U��Q�UV�uW�}�E� �E�P�ER��QPVW�Y�����i��   ���_^��]� ����U��Q�U�E� �E�P�ER�U��Q�MPQR�[�������]� ��U��V�u�~r�FP�*�  ��3��F   �F�F^]� ���U��S�]V�u;�t!W�}j�j V����������;�u��_^[]ËE^[]����������U����Pg3ŉE����M;�tT�PS�XV�p�]��YW�x�X�Y�X�Y�X�Y�X�Q�U��q�q�y�Q�P�p�q�Q�P_�p^�Q[�M�3��e ��]� ���U��j�h��d�    PQV�Pg3�P�E�d�    ��u��v 3��N��j��A�A   P�E��A�EP�����ƋM�d�    Y^��]� �������U��EVP�������4���^]� ����U��V�����~$r�FP��  ��3��F$   �F �ΈF� �Et	V��  ����^]� ������U��j�h��d�    PQV�Pg3�P�E�d�    ��u�� 3��N�(�j��A�A   P�E��A�EP�+����ƋM�d�    Y^��]� �������U��Q�V�u3�j���R�F   �VP�ΉU��V�������^��]� �������������U��j�h4�d�    P��   SVW�Pg3�P�E�d�    3ۉ]��}����   9��   j�v�  �����u3��E�;�t2�M�E�P�Y���P��`����E��E�   ����j P�λ   ������E�   ���t�����`����]��t�����t�}�r�M�Q� �  ���   �M�d�    Y_^[��]�������V���(��~$r�FP���  ��3��F$   �F �F��^�� ��������������U��V���(��~$r�FP��  ��3��F$   �F �ΈF� �Et	V�`�  ����^]� ������U��UV���W�F   �F    �F �x�@��u�+�PR������_��^]� �����U��Q�UV�u3��F�F   �E��F�EPRQ���������^��]� �������������U��j�hh�d�    P��4�Pg3ŉE�SVWP�E�d�    �]�щUЃ��u3��  �B$���t �B4�0�;�s��B$��Q������  �BL����  �z< uP��P�� �������  ����  �   3��E� �]̉M�E؉E��E�   ��s�E��@ �E�    �E؋U�I ���	  �؉]ȅ�t!�ȃ�s�M�;�w�ȃ�s�M؋u��;�v� �U�E؍Mԃ��t�ȃ�s�M؋u��;�r�Y �U�E؋}����  ����t$�ȃ�s�M�;�w�ȃ�s�M؋]�ˋ]�;�v� �U�E؍Mԃ��t��s�E؋U��;�r�� �EЋH<��R�E�P�SV�E�P�E�P�E�P�EЃ�DP�҅���  ���9  �U�E؃��  ����t!�ȃ�s�M�;�w�ȃ�s�M؋}��;�v� �U�E؍Mԃ��t�ȃ�s�M؋}��;�r�Z �U�E؋}�+�tz����   ����t!�ȃ�s�M�;�w�ȃ�s�M؋]��;�v� �U�E؍Mԃ��t��s�E؋U��;�r�� �EЋHLQWjV�" ��;���   �U�E؋M��AA�M�9M�u|�������}� �M�s{j j�S���������]؉]�������u��Q����u�������u��D�����uB�UЋBL�M�PQ��������t�u�M��������'�Mԃ����������M��y����E��M��l�������M�d�    Y_^[�M�3��m ��]� �����������U���SV��F W�~@98u�}u�~< u�]K��]�~L ��   �G�����tw��u�}t�M�VLQSR��" ����uX�NL�E�PQ��! ����uD�V 9:u�N�9�V �FA�Ή�V0+ȃ�A�
�E�M��U�_�H�ND^�     �P�H[��]� �E�x�_3�^��H�H�H[��]� �������������U����EV��~L �MW�}�E��M���   ���v�����t�FL�U�RP�" ����uk��t�NLjWQ��! ����uT�FL�U�RP��  ����u@�M�V �ND�N@9
u�FAPPQ��������E�M��U��H�ND_�     �P�H^��]�  �E�x�_��@    �@    �@    ^��]�  �����������U��QSVW�}���    ��t�E9Fw;Fv� �E�]���G9^w;^v� �]����t;�t�� �G;�tB�VPRS�V����؋F���E���;�t��I ���)������   ;}�u�E_�^^[��]� ��_^[��]� ����S��V�s3�;�t(W�{;�t����������   ;�u�CP��  ��3�_^�C�C�C[����������������SV��3�W��9^Lt������u3��FLP�! ����t3��Έ^H�^A�����^L��}��_�^<�ND^[����U��j�h��d�    P��D�Pg3�P�E�d�    jhH��M��E�   �E�    �E� ������E�P�M��E�    ����hl?�M�Q�E�4�� ��U��j�h��d�    PQVW�Pg3�P�E�d�    ��u��}W�U 3�j��N���GR�A   �QP�U��Q�����ƋM�d�    Y_^��]� �U��EVP�������4���^]� ����U��j�h��d�    P��SVW�Pg3�P�E�d�    j �M��� �=�~ ��}�E�    �]�u+j �M��g� �=�~ u��~@��~��~�M��n� �}�5�~�;ps"�H����u�x t��� ;ps�P�4��3�����uN��t���F�E�WP���������uh\��M�� h�?�M�Q�  �u��Ή5�}�yh��V�`� ���M��E�������� �ƋM�d�    Y_^[��]��������������U��Q�U�E� �E�P�ER�U��Q�MPQR��������]� ��U��j�h�d�    P��   SV�Pg3�P�E�d�    �E3ۉ]�����   9��   j��  �����u�]���t7�M�E�P�|���P��\����E��E�   �5����   �F    �D��3��M�E�   �1��t�����\����]�������t�}�r�U�R��  ���   �M�d�    Y^[��]�U����US�]V�uW�}2��E��M��E��E�PQRWVS�����+�$I�������������    +ȍ�_^[��]��������U��V�uW�};�t*S3ۃ~r�FP��  ���F   �^�^��;�u�[_^]����U��Q�E�V�u3҉j��N��R�A   �QP�U��Q�@�����^��]����������U��j�hQ�d�    P��SVW�Pg3�P�E�d�    �e��u�}3ۉu�]���$    ;}tY�u�u��E�;�tj�S�F   �^W�Έ^��������]��u���ǋu�};�t�]V���R�����;�u�3�SS�I �ƋM�d�    Y_^[��]���������������U��j�h��d�    P��   �Pg3�P�E�d�    �E���A�I#���   �} t	j j �� ��t5h���M������E�P�M��E�    ����h�@�M�Q�E�@�� ��t5h���M��y����U�R�M��E�   �F���h�@�E�P�E�@��h hh���l����A�����l���Q�M��E�   ����h�@�U�R�E�@��- �M�d�    Y��]� �����U��j�h��d�    PQVW�Pg3�P�E�d�    ��u��}W�� 3�j��N�(��GR�A   �QP�U��Q�����ƋM�d�    Y_^��]� �U��EVP�������@���^]� ����U��QS3�V��WSS�^$�^�^�F  �F   �^�^�^ �.���j��  ����;�t6�� ���� j �M������ �C���s@�C�M���� �~$_^[��]�_�^$^[��]���������������U��j�h��d�    PQV�Pg3�P�E�d�    ��u��E�    �����P���  ���M�d�    Y^��]�U��j�h��d�    PQVW�Pg3�P�E�d�    ��u�����~H �E�    t�����~8�E����������t���3c��W�}�  ���N�Z� �M�d�    Y_^��]��U��V���u����Et	V�I�  ����^]� ���������������U��j�h�d�    P��SVW�Pg3�P�E�d�    �E�P�c��P�E�    �����}������E�������t;j �M��Q� �G��v	���sH�G�w����֍M�#��V� ��t
��j���Ћ�E�RP���ҋM�d�    Y_^[��]� ���U��V3�W�}��F�F�F;�u_2�^]� ��I�$	v����PW�;�������    +ύ��F�F_�V�^]� �����������U��j�h@�d�    P��   �Pg3ŉE�SVWP�E�d�    �e��ًC��u3���K+ȸ���������������} �C  �s��+K�������ыM������º"""+Љ�p���;�s�L����;��  ����"""+�;�s3���;�s��j W�����u+s�ȸ������E������P���U������p���+ƍ�RQ���E�    �������p����E�KRPQ�������U��p�������+ƍ��C�MRPQ���o����s�K+θ��������������E��t	V��  ����p�������+ύȋM�S����+эЉK�C�  ��p���R�}�  ��j j �8 ��+M�u��������������¹   ��t����;Esy�}�E��p�������+�����QRP�������K+M��t���P�������C��������+�WP���E�   �����s�[�E��t���R+�SP�`������N�E����+���p�����P���P+�W���7�����p����UQWR�C������t���P�E�VP�������M�d�    Y_^[�M�3��q� ��]� ���������������U��j�h��d�    P��  SVW�Pg3�P�E�d�    �e���u�F��u3���N+ȸ��Q��������ڋ}����  �N��+V���Q��������º�G+�;�s�����8;��g  �����G+�;�s3���;�s��j S�*����U+V�ȸ��Q��������E�i��   3҃��U��U��UR�W�M�P�������E�M�VPQR���E�   �1����E�N�U�i��   E��E�   PQR�������N�V+Ѹ��Q�����������E�������t�VRQ���
����FP��  ���E�i��   i��   ���^�~�F�M�d�    Y_^[��]� �]����u�}�~��i��   �Q�M�W������~ �U�M�i��   i��   �P�V����W�b�  ��j j � +M���Q���������;���   �UR�����軺���E�V��i��   �QRP���E�   ������N��+U�����P���Q���������+�WQ���E��*���^�v�U�����Q+�VR�E�   �z�����������   �E�M�i��   �Q�R�U�P����j j �M �EP��P�������i��   �^S��+�SP���E�   �E�F����M�USQR�F�������P���P�E�WP���������P����E������=����M�d�    Y_^[��]� ���������U��QV��VW��u3��
�F+����ȋ}����  S�^��+�������?+�;�s�}����8;���   �������?+�;�s�E�    �M��ȉM�;�s�U���j Q�Ѽ���]+^�M��Q��W��R�ΉE��&  �E�M�VPQR���&  �V�;�]���EQRP���f&  �F�N+������t	P��  ���U������^[_�F�N^��]� �E��+���;�s]�M���    �M�QSP�ΉU�&  �F��+U�MQ��+�WP���+&  �EF�v�U�MQ+�VR�%  ��[_^��]� �E���    S��+�S�MW�ΉE�%  �USWR�F�h%  �M�EP�E�QP�5%  ��[_^��]� ���������U��Q�M�U�E� �E�P�EQ�MR�UPQR��������]�����U��j�h��d�    P��SVW�Pg3�P�E�d�    j �M��Z� �=�} ��}�E�    �]�u+j �M��7� �=�} u��~@��~��}�M��>� �}�5�}�;ps"�H����u�x t��� ;ps�P�4��3�����uN��t���F�E�WP�l��������uh\��M��o  h�?�M�Q�� �u��Ή5�}�IX��V�0� ���M��E������� �ƋM�d�    Y_^[��]��������������U��V�uW�};�tS�]j�j S���������;�u�[_^]������U��Q�E�MV�uPQV�E�    �3�������^��]����������U��j�h��d�    P��SVW�Pg3�P�E�d�    �e��u�}3ۉu�]���$    ;�vZ�u�u��E�;�t�Ej�S�F   �^P�Έ^�#���O���]��u�ǋu�};�t�]V��������;�u�3�SS� �M�d�    Y_^[��]�U��j�h��d�    PQV�Pg3�P�E�d�    �M��A��P�D
����q����E�    �����F��H�D1����M�d�    Y^��]�������������U��EVWP���@�������B�����Є�t�G<    _^]� �ωw<�W���_^]� �U���   �Pg3ŉE�SV�ًCW�   �u�}��{�u��+ȸ��������������;�vH9{v� �K+K�E�P���������������+�VWP������_^[�M�3��� ��]�| s]9{v�: �K���t����M�;Kv�" �M���M�V��|�����|����������t����M���|���WPQR��t���P��������M�_^3�[�/� ��]�| �������������U��j�h�d�    P��SVW�Pg3�P�E�d�    ��^�F�}��+ȸ��Q����������E�    ;�v59^v�j  �V+V��EP���Q���������+�WSQ���:����PsN9^v�3  �F��M�E;Fv�  �E��E�W�E�P�M�U�������M�P� SQRP�M�Q�������M�E������I����M�d�    Y_^[��]�� �����U��E�UP��Q�MQR�X�����]� �U��j�hH�d�    PSVW�Pg3�P�E�d�    ��3�9^L��   �E�M�UPQR�d� ����;���   ���FH�^A�±���O�N0�N4�G�M�F�F�~ �~$�~L��}Q�ΉFD�^<�Q���P�]��H�������B�����Є�t!�M�^<��S���ƋM�d�    Y_^[��]� �Ή~<�K����M��S���ƋM�d�    Y_^[��]� 3��M�d�    Y_^[��]� �������U���SV��FW�~��+�������u3��#;�v�m� �M���t;�t�[� �]+����U�E�MRjPQ�������~;~v�1� �6�u��}���u� � 3��<�;xw��t�6����3�;~s��� �E�U��x_^�[��]� ���U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U��j�h��d�    P��4�Pg3ŉE�SVWP�E�d�    �e��u�}3ۉủu��E�   �]�]ԉ]��E�;}te�uĉu��E�;�tj�S�E��F   �^P�Έ^����W���E��������ũ�뻋uȋ}�;�t�]V��������;�u�3�SS�� �}�r�M�Q�7�  ���ƋM�d�    Y_^[�M�3��&� ��]�������V�qX���5���V�|��� ��^�����V���HW�13��@u�@(��ȋB0�Ѓ��u�   ��I΅�t�Aǃy( u��j P�E���_��^�U��QV��F��t�M�Q�N�VRQP������VR�w�  ���P�F    �F    �F    �W�  ��^��]����������������U���V��NW��u3���F+����~��+���;�s�E�����~_^��]� ;�v�� �U�RWP�E�P������_^��]� ������������U��VW�y��wX�������V�|��D� ���Et	W裲  ����_^]� ��������U��j�h��d�    P��SVW�Pg3�P�E�d�    �e���u��H�D1΅��(  �I,��t�Q����} ��   ��P�L2����   �MQ����8P��P�E�    ��������M���O����B�L0(�A �8 �E�   t�Q0�: ~� � ���P�҃��u!��H�D1΃��y( u��j P�L�����W���JHu*�E�������H΃y ue��M�d�    Y_^[��]� ��H�L1(�ֿ��딋M��B��H���x( u�����H�Hu�E�������HËu��j j ��� �A���y( u��j P����2��M�d�    Y_^[��]� ��������U��SVW�}���    ��t�E9Fw;Fv�� �E�]���G9^w;^v�d� �]����t;�t�P� �O;�t5�F�E �UR�UR�URQPS�w����V�؋EP�NQRS�������(�^��_^[]� ����U��Q�UV�uW�}�E� �E�P�ER��QPVW��������    +΍�_^��]� ��U��SV�uW�}��+ϸ�$I�����������    +ȋE�ɋ�+�;�t+ƉE��E��V�0�����;�u�_^��[]�����U��j�h��d�    PQV�Pg3�P�E�d�    ��u��E���Q�D(��t�H�l� �E�P�E�    ������F�ƋM�d�    Y^��]� ����U���SV��FW�E�9Fv��� �~�;~v��� �M��QSWP�U�R������_^[��]������������U��j�h7�d�    P��SVW�Pg3�P�E�d�    ���}�3��E�9Et����GX���E��E�   ��Q����G��p���������_j �Ή^(�F,    �?����~( �F0u�F����j P��������F    ��Q���E�   ����B���������CH �CA �M���3��CL��}�C<�KD�ǋM�d�    Y_^[��]� ������U��j�h��d�    P��SVW�Pg3�P�E�d�    ���}�3��E�9Et����GP���E��E�   ��Q����G��p���������_j �Ή^(�F,    �?����~( �F0u�F����j P��������F    ��Q�E�M��PQ���E�   ���������ǋM�d�    Y_^[��]� �U��j�h��d�    P��SVW�Pg3�P�E�d�    �e���u�   S3�V�M��}�~�����}� �}���   �}��~{��H�L1(�A �8 �]�t�Q0�: ~� � ���P�҃��u	]��@�M;�u.^��H�L1(�Q �: t�A0�8 ~	��I ���B���
+���s�M��E�    �}�M� �~ u����J��΅�tA�y( u��j P�����E���Q�D(�E�������t�H��� �ƋM�d�    Y_^[��]� ^�M�ˉM��Q�L2(�'����'����M��@��H���x( u�����H�Hu�E�    �oNËu��?���j j �7� ����������������U��j�h��d�    P��SVW�Pg3�P�E�d�    �e��u3�WV�M܉}��E� �o����}� �}���   ��I�E�P��"I��P�E��������M���E� �H���Mj�W�L�����B�0�A�E���~�����r������I(�A �8 t�Q0�: ~� � ���P�҅�v	���uy�M��E�    �}��@ƀ}� �@    u����I΅�t�Aǃy( u��j P������E܋�J�D(�E�������t�H�6� �ƋM�d�    Y_^[��]ËS���JH�{����MPj�_�����H�L1(�E�O�\����K����M��B��H���x( u�����H�Hu�E�    �:PËu�&���j j �l� �����U��Q�U�E� �E�P�ER�U��Q�MPQR�{�������]� ��U��Q�M�U�E� �E�P�EQ�MR�UPQR�;�������]�����U��QVW�}��;��W  �G�O+ȸ�$I����������Eu�������_��^��]� �NS�^+˸�$I�����������9MwY�GSP�GP�����MQ�N�VRQP�����O+O��$I�������������    +ЋF[��_�N��^��]� ��u3���V+ӉU���$I���U��������9Ew+�G��    +э�SQP�M������F�O�U��PQR�M��t�FPS�������FP��  ���O+O��$I�����������P���q�����t�N�W�GQRP�������F[_��^��]� ������������U��j�h �d�    P��X�Pg3ŉE�SVWP�E�d�    �e��E��E��F�u���u�E���N+ȸ�$I����������E��}����  �^��+N��$I����������¹I�$	+�;�s������M��;��  ����I�$	+�;�s�E�    �M��ʉM�;�s�E���j Q�ܥ���]+^�ȸ�$I��������3���ڋU����E��E�R��    �M�+Í�WQ�Ή]��W����U��E�NRPQ���E�   ������E�ߍ�    +Ӎ��V�EQRP���E�   ������^�N+˸�$I��������������t�VRS���(����FP�/�  ���E���    +ȋE�����    +ωV���V�F�  �]����u��}�~��    +ƍ�Q�M�W�������~(�U���    +ȍ���    +ƍ�RQ�M�����W誥  ��j j �e� +]��$I�����������;���   �M�Q�M������E�N��    +��ۍRQP���E�   �����N+M�U�R��$I�����������+��FWP���E������^�v�U�M�Q+�VR�E�   �!������M��   �M��    +��M��Q���R�U�P�����j j �� �E�P�M�������F��    +��P���P+�W���E�   �E�������M��UQWR�F�����E�P�E�SP�������M��Y����M�d�    Y_^[�M�3��]� ��]� �����������U��j�h[�d�    PQV�Pg3�P�E�d�    ��u��E��F�@   �@    �@ ��E�    ��t0PQ������Q���D��t�    �M�d�    Y^��]� �ƋM�d�    Y^��]� ������������U���SV��^W�~��+ϸ�$I�����������u3��3;�v� � �M���t;�t�� �M+ϸ�$I������������M�U�EQjRP���j����^;^v��� �6W�M��u��]��ܠ���E�M��U�_^��P[��]� �����U���SVW���G��u3���O+ȸ�$I�����������_��+O��$I�����������;�s.�U�E� �M�Q�MR�GPQjS���������__^[��]� 9_v�"� �U�RSP�E�P������_^[��]� ���������������U��j�h��d�    PW�Pg3�P�E�d�    �}�E�E�   ;E,tP��u�� �ML�EP�����E��u�� �E��t#�MQP�y�����J���Dt3��E��E;E,u��}(�UL�r�EP觡  ���}H�E(   �E$    �E r�M4Q胡  ���ǋM�d�    Y_��]���������������U��j�h��d�    P��V�Pg3�P�E�d�    �ML�UL�E� �E�P�ELQRP�� �̍U,�e�RQ�E�   �]������čM�e�QP�E��G����u��V�E�������T�}(r�UR�ՠ  ���}H�E(   �E$    �E r�E4P豠  ���ƋM�d�    Y^��]�������������U���}��t]��]���������������̡�}���   ��}ǀ�   `Y�p   �������������������������������U��E�� t��t3�]ù�}�C �����]ø   ]����j j j jdjdhZ� j���  � ����U��j�hI�d�    P��VW�Pg3�P�E�d�    h�jh ~jH�f�  ���E��E�    ��t����   ���3���}�H�A�U�R�E������Ћ�}�Q�Jj j��E�h�P�у��U�R�M��E�   ��M �0Wj�E��8 ��PVj j�8 ��PhZ� �%J ���M����E���N ��}�H�A�U�R�E������Ѓ��ƋM�d�    Y_^��]��������G �����������U��j�h��d�    PQV�Pg3�P�E�d�    ��u��RG �N�E�    ��������ƋM�d�    Y^��]������������U��j�h��d�    PQV�Pg3�P�E�d�    ��u��N�E�    �������E�������F �M�d�    Y^��]�����������U��V�������Et	V��  ����^]� ����������������x�����������U���EV���x�t	V訝  ����^]� ��������������U��U�BV�uW�}�g��'���F�g��'��������������AzT�M�B�f��&���A�f��&����������u.��!�B�a����!�G�a����������u_�   ^]� ��_3�^]� �������������U��M��t	��Pj��]������������U�����SV�U��Nh+Nd����*���������3�;ÉE�H���   �I����]��E�W�Vh��+Vd����*���������;�r�� �Nh+Nd�~d}�����*���������;�r��� �U��Fd�D�����G�U��C��;]���U��E��U�|�_���^[��]����������U��E��SV��Nh+NdW�}������*���������;�r�� �Fd�[�ЋU���M��Nh+ȸ���*���������;�r�R� �Vd�[�ʋM���Nh�E�+ʸ���*���������;�r�!� �Vd�E��[�D����`�U���M�� ���B�`�� �����^����z_^2�[��]� 3�9]~]�;]tQ;]tL;]tG�Nh+Nd�<�����*���������;�r�� �Vd��ʋM�U�P�E�QRP���A�����u��}C;]|�_^�[��]� ���������V��W����F|3�;�t	P藚  ���FpP�~|���   ���   �|�  �Fd��;�t	P�l�  ���NXQ�~d�~h�~l�W�  �FL��;�t	P�G�  ���V@R�~L�~P�~T�2�  ��_�x�^�������U��j�h��d�    PQV�Pg3�P�E�d�    ��u��N@�E�    ����"  �NX�E��  �Np�E��
  �ƋM�d�    Y^��]���������U��j�h�d�    PQ�Pg3�P�E�d�    h�   胗  ���E��E�    ��t���K����M�d�    Y��]�3��M�d�    Y��]������������U���S�ًKh+Kd����*����W��������]��y  3ɋǺ   ����V���Q���  ���ˋ��E� �����@�����Au3���~'��$    ��@;�|��3���~�O���@I;�|��E����ߍ?�G���   ��M��E���I�M�����   ;؋ȉM�
�E�    �M�A;؉E�
�E�    �E��x;�3�VSWPQ�M��L�������   �}� �E�M������<��E�U�t-�M�E��E�P������M�U��M��MR������M�E��}�P�.�}��}�M�Q�������U�E�P�ωU������M�U�M�R�������E�@;�}����L��@;�|�K��U�������V�ޗ  ��^_[��]� ��U��]�G����������U��M����w3ɍI���R�b�  ����]Ã��3����sލEP�M��E    �� h�;�M�Q�E�h���� �������U��E�M;�t�UV�2�0��;�u�^]��U��E�U+���V�u��    +��~QRQV��� ����^]�U��E�U+�V��W�}��    �49��vQRQW�� ��_��^]� �����������U��V�uW�}�Ƌυ�v�US��H����w�[��_^]� ���V��F��t	P�P�  ���P�F    �F    �F    �0�  ��^������������U���E��P���\$�E�\$�E�$��]� �����������U��VW�����u�� ���t��3ҋE�4@�G����;Bw��t�	�3�;As�_� w��_^]� �������������U��E�U;�t.�MV�1�0�q�p�q�p�q�p�q�p�q�p��;�u�^]����U��M�U�E;�t.V�1�0�q�p�q�p�q�p�q�p�q�p����;�u�^]�U��U�M�E;�t0V�q���p�q���p�q�p�q�p�q�p�q�p;�u�^]���������������U��V��NP+NL����*��������W�}�;�r�M� �VL��ʍʋM�U��@_�^�@�E�]� ���������������U��V��NP+NL����*��������W�}�;�r��� �VL��ʍʋM�U��@_�^�@�E�]� ���������������U����US�]V�uW�}2��E��M��E��E�PQRWVS�����+󸫪�*��������@������ȋ�_^+�[��]�������U��M�U�E;�t2V��t"�1�0�q�p�q�p�q�p�q�p�q�p����;�u�^]�������������U����US�]V�uW�}2��E��M��E��E�PQRWVS�����+󸫪�*����������@��_^[��]����������������U��U��v6�M�EV��t"�1�0�q�p�q�p�q�p�q�p�q�pJ����w�^]���������������U��Q�M�U�E� �E�P�EQ�MR�UPQR�{�������]�����U��Q�UV�uW�}�E� �E�P�ER��QPVW�Y����v����_^��]� ��������U��SVW�}���    ��t�E9Fw;Fv��� �E�]���G9^w;^v�� �]����t;�t�� �G;�t�VPRS�w������F��_^[]� ��������U��S�]V��W�    ��t�E9Fw;Fv�@� �E�}���C9~w;~v�$� �}����t;�t�� �S;�t/�F+�����    ���~QWQR�0� ���E_�^^[]� _^��[]� ����������U��Q�U�E� �E�P�ER�U��Q�MPQR�K�������]� ��U���SV��FW�E�9Fv�|� �~�;~v�m� �M��QSWP�U�R���r���_^[��]������������U���SV�ًCP�s@W�E�9Fv�)� �~��E�;~v�� �M��U�QRWP�E�P�������{h9{d�sXv��� ��M�N�M�;Nv��� �M��U�WRQP�E�P����������   9{|�spv�� �^��M�;^v�� �U�WRSP�E�P���$���_^[��]��������������U��V�������Et	V詏  ����^]� ���������������U��j�hp�d�    P�� SVW�Pg3�P�E�d�    �e���F��u3���V+и���*��������ȋ}���V  �^��+V����*��������º���
+�;�s������8;��  ���軪��
+�;�s�E�    �M��ȉM�;�s�U��j Q�P����U+V�ȸ���*��E���ڃ����P�[��W�MP���E�    �'����M�U�FQRP���t����Uߍ[�ʋN�UPQR���Y����^�N+˸���*������������t	S�D�  ���E�@�E�ȍ�V�ȉV�F�M�d�    Y_^[��]� �EP�	�  ��j j ��� �M��+Ѹ���*���������;ǋE��   ��UԋP�U؋P�U܋P�U��P�@�E�����E�PSQ�ΉU������^�M�Q��+M����*���������+�WS���E�   � ����EF�v�U�M�Q+�VR��������M�d�    Y_^[��]� ��P�MԋH�<�U؋P��M܋H�U��P�S���+�S�M�P�ΉU�E������M�F�ESPQ�R����E�U�R�WP�R������M�d�    Y_^[��]� �����������U��j�h��d�    PQV�Pg3�P�E�d�    ��j蓊  3Ƀ�;�t�0�3���N�N�N�ƋM�d�    Y^��]��������U���SV��^W�~��+ϸ���*���������u3��1;�v��� �M���t;�t��� �M+ϸ���*����������M�U�EQjRP���^����^;^v�� �6W�M��u��]�������E�M��U�_^��P[��]� ���������U���SV��^W��u3���N+˸���*��������ʋ~��+Ӹ���*���������;�s.�U�E� �M�Q�MR�FPQjW�\��������~_^[��]� ;�v��� �U�RWP�E�P������_^[��]� �����U����QP�E+QL��V�U��E�q@����*�����U��E���U��������u,���������Q�Y(�Q�Y0�Q �Y8�M�Q��� ���^��]� �������A������Au���Q���Q����z�Q�A ������Au���Q ���A(������z���Y(����A0������z���Y0����Q8����A�z����M���Q���{���^��]� ����U��E�E��$V3��0W���_�OP+OL����*�����������  S�OX�����G(�g�G0�g�G8�g ��������Au.������Au%�؉u�������Au	�E   �o�   �E   �f������z2��������Au+���E�   ������Au3��E   �5�   �u�+����������E�   ����z3��E   ��u�   �OP+OL����*��OP+OL������򸫪�*���������u�� �GL��vI�M�ȉU��U��؉M�А��E�M��]�� �U��]�R��OX�]������   EE�؃�u͋��   �wp�E9Fv�N� �^��E�;^v�<� �M�U�QRSP�EP������V���&����N+N���������E��[�t�N+N����w��� �F_^��]� _3�^��]� _��^��]� ��%��%��%��%���U��E��}� ]�̡�}�P�BVj j����Ћ�^���������U���}�P�E�RVj P���ҋ�^]� U���}�P�E�RVPj����ҋ�^]� ��}�P�B�����U���}�P���   Vj ��Mj V�Ћ�^]� �����������U���}�P�EPQ�J�у�]� ����U���}�P�EPQ�J�у����@]� ���������������U���}�P�E�RtP�ҋ�}���   P�BX�Ѓ�]� ���U���}�P�E�Rlh#  P�EP��]� ���������������U���}�P�E�RlhF  P�EP��]� ���������������U���}�P�E�RtP�ҋ�}���   �M�R`QP�҃�]� ���������������U���}�P���   ]��������������U���}�P�E���   P�҅�u]� ��}���   P�B�Ѓ�]� ��������U���V�u�W�}�����Dz�F�_����D{:�F����$�:� �G��$�]��*� �E���������D{_�   ^��]�_3�^��]���������U���VW�M��`����E�}��t-��}�Q4P�B�Ѓ��M��u����_3�^��]Ë�R(���}�H0�QW�҃��M��tԋ�R Q�MQ���ҋ��}�P�B �M��Ѓ��t��}�Q0�Jx�E�PW�у��M��.���_��^��]�������U���}�P�B VW�}�����=NIVb��   ��   =TCAbtR=$'  t6=MicM��   ��}�Q���   j hIicM���ЋWP�B����_^]� ��BW����_�   ^]� ��}�Q���   j hdiem���ЋWP�B����_^]� =INIb��   �~ u���B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� ��  _3�^]� =cnys����_3�^]� ������V�������}�H0�Vh�t�҉F���F    ��^�����V��F�����t��}�Q0P�B�Ѓ��F    ^�����̡�}�P0�A���   P�у����������U���}�P0�E�I���   PQ�҃�]� �������������̡�}�I�P0���   Q�Ѓ���������̡�}�P0�A���   j j j j j j j j j4P�у�(������̡�}�P0�A���   j j j j j j j j j;P�у�(�������U���}�P0�E�IPQ���   �у�]� ��������������U����E V��P�M��;�����}�E�Q�R4Ph8kds�M��ҡ�}�E     �H0���   �U R�U�E�P�Ej R�UP�ER�UP�FRj2P�ыu ��(�M��������^��]� ��������������̡�}�I�P0���   Q�Ѓ����������U��V��F��u^]� ��}�Q0�M ���   j j j j j Q�Mj QjP�ҡ�}�H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uË�}�Q0P�B�Ѓ������̋A��u� ��}�Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5�}�v0Q�MQP���   R�U�R�Ћu�    �F    ��}���   j P�BV�Ћ�}���   �
�E�P�у�$��^��]� �������U���}�P0�E�I�RPQ�҃�]� �U��A��t)��}�Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5�}�v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5�}�v0QP���   R�Ѓ�^]� �����������U��Q��u3�]� �E�H� V�5�}�v0Q�MQPR�V\�҃�^]� ����������U��y u3�]� V�u�W�}�؉��ډ��}�P4�A�JhWVP�ы�ډ����ى_^]� �����U��A��u]� ��}�Q4�M�RhQ�MQP�҃�]� ����U��A��u]� ��}�Q4�M�RpQ�MQP�҃�]� ����U��y u3�]� V�u�W�}�؉��ډ��}�P4�A�JpWVP�ы�ډ����ى_^]� �����U���$VW��htniv�M��	�����}�P�E�R4Phulav�M��ҡ�}�P�B4hgnlfhtmrf�M��Ћ�}�E�Q�R4Phinim�M��ҡ�}�P�E�R4Phixam�M��ҡ�}�P�E�R4Phpets�M��ҡ�}�P�E�R4Phsirt�M��ҋE �}$=  �u�����t.��}�QP�B4h2nim�M��Ћ�}�Q�B4Wh2xam�M��ЋU�M�QR�E�P���K�����}���   P�B8�Ћ�}���   �
���E�P�у��M��(���_��^��]�  ��������������U���$V��htlfv�M������E��}�P�B,���$hulav�M��Ћ�}�E,�Q�R4Phtmrf�M����E��}�P�B,���$hinim�M����E��}�Q�B,���$hixam�M����E$��}�Q�B,���$hpets�M��Ћ�}�ED�Q�R4Phsirt�M��������E0��������Dzw���]8����Dzm�؋�}�E@�Q�R4Phdauq�M��ҋM�E�PQ�U�R���������}���   P�B8�Ћ�}���   �
���E�P�у��M��������^��]�@ �١�}�P�B,���$h2nim�M����E8��}�Q�B,���$h2xam�M����V�����U���$V��hgnrs�M��*����E��}�E��E�   �Q���   �E�Pj�M��ҡ�}���   ��U�R�ЋM��}�M����E�   �B���   �M�Qj�M��ҡ�}���   ��U�R�ЋU���M�QR�E�P���������}���   P�B8�Ћ�}���   �
���E�P�у��M�������^��]� �U���$V��hCITb�M��J�����}�P�E�R8PhCITb�M��ҡ�}�P�E�R4Phsirt�M��ҡ�}�P�E�R4Phulav�M��ҋM�E�PQ�U�R��������}���   P�B8�Ћ�}���   �
���E�P�у��M��������^��]� U��E��Vj ��P�M�Q�M�uY  �UPR���)������}�H�A�U�R�Ѓ���^��]� ����������U��E,��UPj ���T$�$htemf�E$�� �\$�E�\$�E�\$�E�$R�O���]�( �����������U��E,��Pj ���T$�U�$hrgdf�E$�� �������������\$�E�����\$�M���\$�E�$R�����]�( ���U��E,��Pj ���T$�U�$htcpf�E$�� ��������\$�E���\$�}�\$�E�$R����]�( ���������������U��Q��u3�]� �E�E�H� V�5�}�v0Q�M Q�M���\$�E�$QPR�V(�҃�$^]� ������U��Q��u3�]� �E�H� V�5�}�v0Q�MQPR�V,�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5�}�v0Q�MQPR�V,�҃�^]� ����������U��Q��u3�]� �E�H� V�5�}�v0Q�MQPR�V0�҃�^]� ����������U��SVW���W��t$�E�H�5�}�^0� �uQVP�C0R�Ѓ���u	_^3�[]� �W��t��E�H� ��}�[0Q�NQPR�S0�҃���t̋W��tŋE�H� �=�}�0Q��VP�G0R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5�}�v0Q�MQ�MQPR�V<�҃�^]� ������U��QV3�W��u3��,�E�H� �5�}�v0Q�MQPR�V,��3Ƀ�9M�������}�M�B�P0VQ�M�ҋ�_^]� ����U��AV��u3��"�M�Q�	�5�}�v0R�URQP�F,�Ѓ�����}�Q�E�M�R4PQ�M�ҋ�^]� ���������������U��A��V��u3��"�M�Q�	�5�}�v0R�U�RQP�F0�Ѓ�����}�E��Q�E�M�R,���$P�ҋ�^��]� �����U�����V���U��V�U��]�W��t$�E�H� �=�}�0Q�M�QPR�W0�҃���u
_3�^��]� �V��t�E�H� �=�}�0Q�M�QPR�W0�҃���tˋV��tċE�H� �5�}�v0Q�M�QPR�V0�҃���t���}�P�M�RH�E�PQ�M��_�   ^��]� �����������U��� ��A�U�V�U�W�]���u3��&�M�Q�	�5�}�v0R�U�R�U�RQP�F<�Ѓ����E�}���t��}�Q�RH�M�QP���ҋE���t��}�E��Q���$P�B,����_��^��]� U���}�P�E���   Vj ��MP�ҋM$�U Q�MR�Uj Q�MR�UQPR���o���^]�  ����������U���}��P�E���   V���$��MP���E8�E@�M,�Uj P���\$�E0�$Q�E$�� �\$���E�\$�E�\$�$R�K���^]�< ������U���}��P�E���   V���$��MP����Ej j ���T$���$htemf�E$�� �\$�E�\$�E�\$�$P�����^]�$ �����������U���}��P�E���   V���$��MP���E$�Ej �� �\$���E�\$�E�\$�$P�C���^]�$ ��������������U���}��P�E���   V���$��MP����j j ���T$�E�$htcpf�E$�� ����������\$�E���\$�}�\$�$P����^]�$ ���������������U���}�� V��H�A�U�R�ЋM�E��Qj �U�RP�M�Q�M�����UPR���������}�H�A�U�R�Ћ�}�Q�J�E�P�у���^��]� ������������U���dV��M��_O  ��}�Q���   P�EP�M�Q�M��P�M���O  �M��!P  j j �E�P�M���P  �MPQ��������}���B�P�M�Q�҃��M���O  �M���O  ��^��]� �����U���P��EV�]���W�}����t��}�Q���$P���   �����]����}�U��UЍE��]ȋQ�M���   PQ�E�P���ҋ�M��P�U�H�M�P�U�H�M��P�F�U��u_^��]� �M�E�Q�	�5�}�v0R�U R���\$�U��E��$RQP�F(�Ѓ�$_^��]� ���������������U���0�E�M���u��}�H���   �҅�u��]� SVW���<~  ��htlfv�MЉu�����E�}��}�X�U�����$��� �]��G�$��� �}�S,�M��$hulav�ҡ�}�P�B4hmrffhtmrf�M��Ћ}���}�M�Y���$�� �]��G�$�w� �}�S,�M��$hinim�ҋ}���}�M�X���$�I� �]��G�$�;� �}�S,�M��$hixam�����}�P�B,���$hpets�M��Ћ�}�Q�B4j hdauq�M��Ћ�}�Q�B4Vhspff�M��Ћ�}�E �Q�R4Phsirt�M��ҋM�E�PQ�M��U�R�n�����}���   P�B8�Ћ�}���   �
���E�P�у��M��K���_��^[��]� U��E��V���u��}�H���   �҅�u^��]� ���n|  �E�F��u3��"�M�Q�	�5�}�v0R�U�RQP�F0�Ѓ����E������M������\$�M��$�|  ��M��P�Q�P�Q�@�A��^��]� ����������U���0���}�]�V���M�]�P���   �E�PQ�M�E�P�ҋ�P�M��Hj �U�P�E P�M��MQ�M�U��UR�U�E�PQR������^��]� ���������������U�����UV�]���E�P�]��ERP������}�Q�M�R@���E�PQ�M�ҋ�^��]� ����������U��A��u]� �M�Q�	V�5�}�v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� ��}�Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� ��}�Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U���}�P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� ��}�Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj>P�ҋE���(��]� ������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5�}�v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M�� �MQ�U�R�M��X ��tm�}��E��tN��}���   P�BH�ЋM��I����tQ�W�7��}�[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M��� ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5�}�v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� ��}�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� ��}�Q0�M�RDQ�MQ�MQP�҃�]� U��A��u]� ��}�Q0�M�RHQ�MQ�MQ�MQ�MQ�MQP�҃�]� ���̋A��uË�}�Q0P�BX�Ѓ�������U��A��u]� ��}�Q0�M�RLQ�MQP�҃�]� ����U��A��u]� ��}�Q0�M�RP��   �QP�҃�]� ��U��A��u]� ��}�Q0�M�RPQP�҃�]� ��������U��A��u]� ��}�Q0�M�RTQ�MQ�MQ�MQP�҃�]� ������������U���}V�u�VW���H4�R�ЋE�F    �~�H� ��}�R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� ��}�Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I��}�R0P�EPQ���   �у�]� ������̡�}�I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u��}� ��}�R0�I�R@V�uVP�EPQ�҃�^]� �����������U���}�P0�E�I�RdP�EP�EP�EP�EPQ�҃�]� �U���}�P0�E�I�RpP�EP�EP�EP�EPQ�҃�]� �U��E�P� V�5�}�v0R�UR�UR�UR�URP�A�NhP�у�^]� ��������U��E� ��}�R0j j j j j j j P�A���   jP�у�(]� �����������U��E� ��}�R0j j j j j jj P�A���   jP�у�(]� �����������U��E� ��}�R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M������E�H� ��}�R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R������M��������^��]� ����������U��E�P� V�5�}�v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5�}�v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5�}�v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5�}�v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U���}�P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U���}�UVj j j j j R��H0�E�Vj P���   jR�Ћ�}�Q0�E�N�RtPQ�҃�0^]� ��U���}�P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡�}�P0�A���   j j j j j j j j jP�у�(�������U���}�P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡�}�P0�A���   j j j j j j j j j(P�у�(�������U���}�P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U���}�P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡�}�P0�A���   j j j j j j j j jP�у�(������̡�}�P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}�M���t��}�P���   j j���Љ�u��t��}�Q���   j j���Љ��}�Q0�E��H�R`VWQ�҃�_^[��]� �U���}�P0�E�I���   P�EP�EPQ�҃�]� �����̡�}�P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V�������}�H0�Vh�t�҉F3��F�F�����F   ��^�������V��F�����t��}�Q0P�B�Ѓ��F    ^������U��E�UVj ��MP�EQ3�9MR��Pj �F    ��
Q��������t�~ t
�   ^]� 3�^]� �U��E�A�I��u3�]� ��}�B0Q�H�у�]� ����U���}�P�B S�]V�����=ckhc��   ��   =cksate=TCAb��   ��}�Q���   Wj hdiem���Ћ���BSW���F   �Ѓ~ ��t��t��u3Ƀ���Q���C���_^��[]� �~ tK��B����^[]� �~ t6��������t+�F    ^�   []� =atnit�MQS���/���^[]� ^3�[]� �U��V��~ ��   W�}����   �$���E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN��}�M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W�h�  ���F    _^]� D�R�`�n�|�������������U��V��~ �  �E W�}�E����   �$�p����]������   �   ���]����A��   �   ���]����A��   �r���]������   �`�E������A��uN��������   �C�E��������u1������A{{�*�E���������E������A�����]����DzU����ء�}�U�H0�F���   j j j j j j j RjP���E �U(��(R���\$�E�$W��  ���F    _^]�$ �I j��������դ����������������U���E �E�Uj���\$�E�\$�E�$PR�w���]�  ���U���E �E�Uj���\$�E�\$�E�$PR�G���]�  ���U���E �E�Uj���\$�E�\$�E�$PR����]�  ��̋�3�� ,��H�H�H�������������VW��3��,�9~u��}�H4�V�R�Ѓ��~�~_^����U���}�P4�E�I�RtPQ�҃�]� �U��U��t3�A��}�I0R���   P�ҋ�}�Q0�M���   QP�҃�]� ��}�P0�E�I�R|PQ�҃�]� ������̡�}�P4�A�JP�у������������̡�}�P4�A�JP�у������������̡�}�P4�A�JP�у������������̡�}�P4�A�J|P�у������������̡�}�P4�A���   P�у����������U���}�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U���}�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U���}�P4�E�I�R PQ�҃�]� �U���}�P4�E�I�R$PQ�҃�]� �U���}�P0�E�I���   P�EP�EP�EPQ�҃�]� ��U���}�P4�E�I���   PQ�҃�]� ��������������U���}�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U���}�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U���}�P4�E�I�R(PQ�҃�]� �U���}�P4�E�I�R,P�EP�EPQ�҃�]� ���������U���}�P4�E�I�R0P�EPQ�҃�]� ������������̡�}�P4�A�J4P��Y��������������U����UV��EP�M�Q�NR�E�    �E�    ������}�H4�V�AR�Ћ�}�Q0�Rhj �M�Q�M�Q�M�Q�M�QP�F�HQ�҃� �} ^t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ��������������U���}�P4�E�I�R8PQ�҃�]� �U���}�P4�E�I�R<PQ�҃�]� �U���}�P4�E�I���   P�EPQ�҃�]� ���������̡�}�P4�A�J@P�у�������������U���}�P4�E�I�RDP�EPQ�҃�]� �������������U���}�P4�E�I�RHP�EPQ�҃�]� �������������U���}�P4�E�I�RLP�EPQ�҃�]� �������������U���}�P4�E�I�RPP�EPQ�҃�]� �������������U���}SV�uW�����   �QV�҃�����   ��}���   �]�QS�҃�S��uA��}���   �Q@�ҋء�}���   �Q@V�ҋ�}�Q4�JPSP�GP�у�_^[]� ��}���   �H�у���uD��}���   �H8S�ы�}�؋��   �H@V�ы�}�J4�WSP�AHR�Ѓ�_^[]� hX�h}  ��   ��}���   �BV�Ѓ�����   ��}���   �]�BS�Ѓ�S��uC��}���   �B@�Ћ�}���   �؋B8V�Ћ�}�Q4�JLSP�GP�у�_^[]� ��}���   �H�у���uD��}���   �H8S�ы�}�؋��   �H8V�ы�}�J4�WSP�ADR�Ѓ�_^[]� hX�h�  �
hX�h�  ��}�Q��0  �Ѓ�_^[]� �U���}�P4�E�I��  P�EP�EP�EPQ�҃�]� ��U���}�P4�E,P�E(P�E$P�E �IP�E�RTP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U���}�P4�E�I�RXP�EP�EP�EPQ�҃�]� ����̡�}�P4�A�J`P��Y�������������̡�}�P4�A�JdP�у�������������U���}�P4�E�I��   P�EP�EP�EPQ�҃�]� ��U���}�P4�E�I�R\P�EP�EP�EP�EP�EPQ�҃�]� �������������U���}�P4�E�I�RhP�EPQ�҃�]� �������������U��V�uW��t��؉�}��t��ډ��}�P4�A�JhWVP�у���t��ډ��t��ى_^]� �U��V�uW��t��؉�}��t��ډ��}�P4�A�JpWVP�у���t��ډ��t��ى_^]� �U���}�P4�E�I�RpP�EPQ�҃�]� �������������U���,V��~ ��   ��}�V�H4�AR�Ѓ} t ��}�Q0�RlP�F�HQ�҃�^��]� ��hARDb�MԉE��E�    �|���P�M�Q�N�U�R������}���   ��U�R�Ѓ��M�����^��]� ������U���}�P4�E�I�RlPQ�҃��   ]� ������������U���}�E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U���}�P4�E�I���   P�EP�EPQ�҃�]� �����̡�}�P4�A���   P�у���������̸   ����������̸   �����������U���}V��H4�V�A$h�  R�Ћ�}�Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U���}�P4�E�I�RxP�EP�EP�EPQ�҃�]� �����U���}�P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}�M���t��}�P���   j j���Љ�u��t��}�Q���   j j���Љ��}�Q4�E��H�RpVWQ�҃�_^[��]� �U��Q��}�P�B SVW�}���3���=INIb�/  �  =SACbvt+=$'  t
=MicM�  ��B$W����_�   ^��[��]� ��R3��E��E�EP�M�Q���҅�t��}�U�H4�E�R�VP�AR�Ѓ�_�   ^��[��]� =ARDb�  ��}�Q���   j j���Ћ�}�Qj �؋��   j���Ћ�}�Qj �E����   j���Ћ�}�Qj �E���   j���ЋM���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>���Y���P���1���P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� ��}�Q���   j hIicM���ЋWP�B ����_^[��]� �������������U���}�P4�E�I�RTh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M��Z�����}�Q4�JlP�FP�у��M��|���^��]��������V�������}�H0�Vh�t�҉F���F    ����F   ��^��������V��F�����t��}�Q0P�B�Ѓ��F    ^������U���}�P�B VW�}�����=cksat`=ckhct�MQW��譾��_^]� �Nj j j j j j �F   ��}�B0���   j j j Q�҃�(��t'_�F    �   ^]� �~ t��P����_^]� _3�^]� ���U���}�H���  ]��������������U���}�H0���   ]��������������U���}�H0�U�E��VWRP���   �U�R�Ћ�}�Q�u���BV�Ћ�}�Q�BVW�Ћ�}�Q�J�E�P�у�_��^��]������������U���}�H0���   ]��������������U���}�H0���   ]��������������U��Ej0P�rj  ��]��������������U��Ej0P�R�  ��P�Ij  ��]�����U��E�M��j0PQ�U�R�W�  ��P�j  ��}�H�A�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P��  ��P��i  ��}�Q�J�E�P�у���]��U��Ej$P�i  3Ƀ�������]����U��Ej$P��  ��P�i  3Ƀ�������]�����������U��E�M��Vj$PQ�U�R��  ��P�Mi  ��}3Ƀ��B�P����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P��  ��P��h  ��}3Ƀ��B�P����M�Q�҃���^��]����U���}�H�U�E���   RPj �у�]���������������U���}�H�U�ER�UP���   Rj �Ѓ�]�����������U���}�P4�E�I�R,P�EP�EPQ�҃�]� ���������U���}�P4�E�I�R0P�EPQ�҃�]� ������������̡�}�P4�A�J4P��Y��������������U��U��V��EP�M�QR���d�����}�H0�E�P� R�U�R�U�R�U�R�U�R�VP�AhR�Ѓ��} ^t(�} t(�E�M�;�~<�U��;�}3�E�M�;�~)�U���} u�E�M�;�~�U��;�}�   ��]� 3���]� �����������U��ESVW�؅�u�Y��}�P�}���   j hdiuM���Ћ���tK;3u	_^3�[]� ��}�Q���   j hIicM����;�u��}�Q���   j h1icM���Шu��3_^�   []� �����U���}�P�BT��(V�uhfnic���Ѕ�t��}�Q�ȋ��   j
�Ѕ���   ��}�Q�RPhfnic�E�P����P�M������M��7����u�E�P���9����M��!�����}�Q�B ���Ѓ��t��}�Q�B ���Ѕ�u��}�Q�B$hfnic���Ћ�}�E�Q�R8Pj
����^��]���������U���}�P0�E�IP�EP�EP�EPQ���   �у�]� ��U���}�P0�E�IV�p� ���   V�uj j j V�uVj Pj=Q�҃�(^]� ����U���}�P0�E�IV�p� ���   V�uV�uj j j�Vj Pj=Q�҃�(^]� ���̡�}�I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V�������}�H0�WVh�t�ҋ}�F�E�F    �F   ����F��}�Q���   ��j hmyal���ЉF��t��t�F    ��}�Q���   j
hhfed���ЉF_��^]� �����������U���}�P�B VW�}�����=ytsdt�MQW������_^]� ��}�B0�N���   Q�ҋ�P������_�   ^]� ��3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ��������������������̸������������U���E�Y(]� ���U���(V���P(�M�Q���ҋN��t&��}�R0j j j j j j P���   j jQ�Ѓ�(��}�Q�J�E�P�ы�}�B�P�M�Q�ҋF����t ��}�Q0�RHj �M�Qj jj?j P�҃���}�H�A�U�WR�Ћ�}�Q�J�E�P�ыF����u3��;��}�E�    �J0�U�Rj j j h  
 j�U�Rh�  jP���   �Ћ}���(��}�Q�J�E�P�у���_u3�^��]Ë�}�B�P�M�Q�ҋF����t ��}�Q0�RHj �M�Qj j j8j P�҃���}�H�A�U�R�ЋF����t��}�Q0jP�BP�Ѓ���}�Q�J�E�P�у��M�����Ph   h  K j;�U�Rh	��h�  ��跶����}�H�A�U�R�Ѓ��M������F��t��}�Q0P�BX�Ѓ��F��t��}�Q0P�BX�Ѓ��F��t'��}�Q0j j j j j jj j jP���   �Ѓ�(j�v$�Q`  ���   ^��]�����U���SV��W�~j���Y�  ��V�^(3ۉ^4�^8�^<��}�H0�Ah�   R�Ћ�}�Q�J�E�P�ы�}�B�PSj��M�h(�Q�҃�SS�E�P�M�Q���E��  �]��i�����}�B�P�M�Q�҃�Sj����  _^[��]���̍A�������������U��VW��~4 tA�I ��}�H��0  hX�hj  ��j
�/i  ��}�HP�V �AR�Ѓ���uQ9F4u�}�QP�Bh�~0���Ѓ~4 t;��}�Q��0  hX�h�  �Ћ�}�QP�Bl�������m���_3�^]� �M�U�N8�V4��}�PP�Bl�~0���Ѓ~4 t%j
�h  ��}�QP�F �JP�у���u�9F4uۋ�}�BP�PhS���ҋ^<�F<    ��}�PP�Bl���Ћ�[_^]� ��U���}�P�B ��@VW�}�����=MicMtI=fnic��   j�M��8����uP���}����M��e�����}�Q�B4jj����_�   ^��]� ��}�Q���   j hIicM����=�����   htats�M��ҭ����}�Q�B0j j�M��ЍM�Q�U�R�E�P���E��  �E�    �̴����}���   �
�E�P�у��M�轭���F�F   ��t��}�J0�QP�҃��EPW���a���_^��]� ���������U��E��V��t3�^]� j�N�A�  j�
]  �F    �v����t��}�H0�QV�҃��   ^]� ��������������j�����  j�\  ��3�����������U��E3�h�����h  ���P�Ej BR�Uj PR�u���]� �U��Q�Q��u3���]� �E�H� V�5�}Q�M�Q�E�    �v0PR�V8�ҋ�����t@�E���t9��}�Q�M�RQP�ҋE�����t��}�QW��P�B��W��3  ��_��^��]� ������U���}��V��H�A�U�R�ЋU���M�QR���D�������u��}�H�A�U�R�Ѓ�3�^��]� �M�Q�M��  ��}�B�P�M�Q�҃���^��]� �������U���}��V��H�A�U�R�ЋU���M�QR��������M���}�P�R8�E�PQ�M�ҡ�}�H�A�U�R�Ѓ���^��]� �������������U���V��M��/  �M�E�PQ���������}���B�U�@<�M�Q�MR�ЍM���  ��^��]� ����U���}�P�E���   Vj ��MP��h���h  �j j jj P�EP���c���^]� ��������������U���}V�uW�����   �QV�҃�V��u,��}���   �Q@�ҋ�}�Q4�J P�GP�у�_^]� ��}���   �H�у���u.��}���   �H8V�ы�}�J4�WP�A$R�Ѓ�_^]� ��}�Q��0  hX�h	  �Ѓ�_^]� �����U���4��}�H�QSVW�}W�ҡ�}�P�u���   ��3�SS�Ή]�Ћ�}�QS�E����   j���Ћ�;��L  �d$ �} ~l��}�Q�J�E�P�ы�}�B�Pj j��M�h,�Q�ҡ�}�P�B<�����Ћ�}�Q�RLj�j��M�QP���ҡ�}�H�A�U�R�Ѓ���}�Q0�E����   VP�M�Q�ҋ��}�H�A�U�R�Ћ�}�Q�J�E�PV�ы�}�B�P�M�Q�ҡ�}�P�B<�����Ћ�}�Q�RLj�j��M�QP���ҡ�}�H�A�U�R�Ћ�}�Q�u���   �E��j ��
S���Ћ�}�Q���   �E�j �CP���ҋ����������_^[��]����������������U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj AQj R�UR��荱��^]� ��������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR�O���^]� ����������U��E�E43҃8��R�U<R�U(���\$�E,�$R�E �� �\$�E�\$�E�\$�@�E�$P�B���]�8 ��������������U��E�@3҃8��E��Rj ���T$�$htemf�E �� �\$�E�\$�E�\$�$P����]�  ���U��E�E 3҃8��R�� �\$�E�\$�E�\$�@�E�$P�j���]�  ������U��E�@3҃8��E��Rj ���T$�$htcpf�E �� ��������\$�E���\$�}�\$�$P�K���]�  �������U��E3҃8��R�UR�UR�UR�UP�EPR����]� U��E3҃8V�u��V��RP�EP�_���^]� ����������U��Q��u3�]� �E�E�H� V�5�}�v0Q�M Q�M���\$���E�$QPR�V(�҃�$^]� ���U���}�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U���}�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U���}��P�E���   V���$��MP�ҋ���u�^�    ^]� ��u�^����D{�   ^]� ��^]� ������U���0���}�U�V�U���M�]�P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�Q�P�Q�P�@�Q�A����  ^��]� ��������U��� ���}�]�V���M�]��P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�@�Q�A����  ^��]� �����U���VW�}�M�;}us��}�P�u���   j htsem���Ѕ�uS��}�QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E��'�����t�E�M�P�w  _�   ^��]� _3�^��]� U���VW�}�M�;}us��}�P�u���   j htsem���Ѕ�uS��}�QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E�������t�E�M�P��  _�   ^��]� _3�^��]� U���SVW�}��;}uz��}�P�u���   j htsem���Ѕ�uZ��}�QP���   hrdem���Ѕ�u=��M�Q�]��M�U�R�}��E�蕲����t�E������$�  _^�   [��]� _^3�[��]� ��������U���4�ESW�}�M�;�t;Et	;E��   ��}�P�]���   j htsem���Ѕ���   ��}�QP���   hrdem���Ѕ�uj�M��U�U܉E��UԉE��]̉E�M�E�P�M�Q�M�U�U�R�E�P�}�������t+�E̋M�������E��X�E��X��  �   _[��]� _3�[��]� ��������U���SVW�}��;}��   ��}�P�u���   j htsem���Ѕ�uj��}�QP���   hrdem���Ѕ�uM��U�M��]���Q�M�]��E�R�E�P�}��x�����t%�E��������E��X�  �   _^[��]� _^3�[��]� ���̋A���X(Q�ȋB$��j j h�����R  ���������������U���}��0VW���H�A�U�R�Ћ�}�Q�J�E�P�ыE���U�RP�M�Q�M�,>����}�J�U�RP�A�Ћ�}�Q�J�E�P�ы�}�B�P�M�Q�ҡ�}�H�Q��V�ҡ�}�H�A�U�VR�Ѓ�����  ��}�Q�J�E�P�у�_^��]� ������������U���SVW�}��;}��   ��}�P�u���   j htsem���Ѕ�ue��}�QP���   hrdem���Ѕ�uH��}�Q�J�E�P�ыM���U�R�E�P�}��E�    �-�����u ��}�Q�J�E�P�у�3�_^[��]� ���U��R�k<�����  ��}�H�A�U�R�Ѓ�_^�   [��]� ��U��V�u���  ��^]� �����������U���L��}SV��H�A�U�R�Ћ�}�Q�J3�Sj��E�h0�P���F(�����S�U�SR�E��  �]�� P�E�P�S����P�M�Q�������P�U�R���b�����}�H�A�U�R�Ћ�}�Q�J�E�P�ы�}�B�P�M�Q�҃�htats�M��}�����}�P�B0jj�M����F(��}�Q�B,���$j�M��ЍM�Q�U�R�E�P���E��  �]��`�����}���   �
�E�P�у�9^4t^��}�BP�PhW�~0���ҋF4;�t�N8Q�Ѓ��F<�^8�^4���}�B��0  hX�h�  �у���}�BP�Pl����_�M�����^[��]� ������U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�E�Y����D{�   ]� �����������U�����u�E�    �Y�E�Y�E�Y]� ��u-�E�Y����Dz�E�Y����Dz�E�Y����D{�   ]� �����U��V�����u#�E�M�U�F�E�N�V�    �F^]� ��u�MQ�VR菝������t�   ^]� �������������U��V��~ �,�u��}�H4�V�R�Ѓ��E�F    �F    t	V�#  ����^]� �������U��V��F�����t��}�Q0P�B�Ѓ��E�F    t	V�"  ����^]� ��������������U���V��3ɍF��H�������}�M��M����   �RQ�M�QP�ҡ�}���   ��U�R�Ѓ���^��]��������������U��V�����u �    ��}�H�A���UVR�Ѓ��#��u��}�Q�Rx�EP�N�҅�t�   ��}�H�A�UR�Ѓ�^]� �������U���}�P�EP�EP�EPQ�J�у�]� �����������̡�}V��H�QV�ҡ�}�H$�QDV�҃���^�����������U���}V��H�QV�ҡ�}�H$�QDV�ҡ�}�U�H$�AdRV�Ѓ���^]� ��U���}V��H�QV�ҡ�}�H$�QDV�ҡ�}�U�H$�ARV�Ѓ���^]� ��U���}V��H�QV�ҡ�}�H$�QDV�ҡ�}�H$�U�ALVR�Ѓ���^]� �̡�}V��H$�QHV�ҡ�}�H�QV�҃�^�������������U���}�P$�EPQ�JL�у�]� ����U���}�P$�R]�����������������U���}�P$�Rl]����������������̡�}�P$�Bp����̡�}�P$�BQ�Ѓ����������������U���}�P$��VWQ�J�E�P�ы�}�u���B�HV�ы�}�B�HVW�ы�}�B�P�M�Q�҃�_��^��]� ���U���}�P$�EPQ�J�у�]� ����U���}�P$��VWQ�J �E�P�ы�}�u���B�HV�ы�}�B$�HDV�ы�}�B$�HLVW�ы�}�B$�PH�M�Q�ҡ�}�H�A�U�R�Ѓ� _��^��]� ���U���}�P$��VWQ�J$�E�P�ы�}�u���B�HV�ы�}�B$�HDV�ы�}�B$�HLVW�ы�}�B$�PH�M�Q�ҡ�}�H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e�����}�Q$�JH�E�P�ы�}�B�P�M�Q�҃���^��]� ����̡�}�P$�B(Q��Yá�}�P$�BhQ��Y�U���}�P$�EPQ�J,�у�]� ����U���}�P$�EPQ�J0�у�]� ����U���}�P$�EPQ�J4�у�]� ����U���}�P$�EPQ�J8�у�]� ����U���}�UV��H$�ALVR�Ѓ���^]� ��������������U���}�H�QV�uV�ҡ�}�H$�QDV�ҡ�}�H$�U�ALVR�Ћ�}�E�Q$�J@PV�у���^]�U���}�UV��H$�A@RV�Ѓ���^]� ��������������U���}�P$�EPQ�J<�у�]� ����U���}�P$�EPQ�J<�у����@]� ���������������U���}�P$�EP�EPQ�JP�у�]� U���}�P$�EPQ�JT�у�]� ���̡�}�H$�QX�����U���}�H$�A\]�����������������U���}�P$�EP�EP�EPQ�J`�у�]� �����������̡�}�H(�������U���}�H(�AV�u�R�Ѓ��    ^]��������������U���}�P(�R]����������������̡�}�P(�B�����U���}�P(�R]�����������������U���}�P(�R]�����������������U���}�P(�R ]�����������������U���}�P(�E�RjP�EP��]� ��U���}�P(�E�R$P�EP�EP��]� ��}�P(�B(����̡�}�P(�B,����̡�}�P(�B0�����U���}�P(�R4]�����������������U���}�P(�RX]�����������������U���}�P(�R\]�����������������U���}�P(�R`]�����������������U���}�P(�Rd]�����������������U���}�P(�Rh]�����������������U���}�P(�Rx]�����������������U���}�P(�Rl]�����������������U���}�P(�Rt]�����������������U���}�P(�Rp]�����������������U�����}�E�    �E�    �P(�RhV�E�P���҅���   �E���uG��}�H�A�U�R�Ћ�}�Q�E�RP�M�Q�ҡ�}�H�A�U�R�Ѓ��   ^��]� ��}�Qh8�h8  P���   �Ћ�}���E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�F  ��3�^��]� �M��U�j IQ�MR�����E�P�  ���   ^��]� ���������������U���}��V��H�A�U�R�Ѓ��M�Q������^��u��}�B�P�M�Q�҃�3���]� ��}�H$�E�I�U�RP�ы�}�B�P�M�Q�҃��   ��]� �U��Q��}�P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U���}�P(�R8]�����������������U���}�P(�R<]�����������������U���}�P(�R@]�����������������U���}�P(�RD]�����������������U���}�P(�RH]�����������������U���}�P(�E�R|P�EP��]� ����U���}�P(�RL]�����������������U���}�E�P(�BT���$��]� ���U���}�E�P(�BPQ�$��]� ����̡�}�H(�Q�����U���}�H(�AV�u�R�Ѓ��    ^]��������������U���}�P(���   ]��������������U���}�H(�A]����������������̡�}�H,�Q,����̡�}�P,�B4�����U���}�H,�A0V�u�R�Ѓ��    ^]�������������̡�}�P,�B8�����U���}�P,�R<��VW�E�P�ҋu����}�H�QV�ҡ�}�H$�QDV�ҡ�}�H$�QLVW�ҡ�}�H$�AH�U�R�Ћ�}�Q�J�E�P�у�_��^��]� �������U���}�P,�E�R@��VWP�E�P�ҋu����}�H�QV�ҡ�}�H�QVW�ҡ�}�H�A�U�R�Ѓ�_��^��]� ��̡�}�H,�j j �҃��������������U���}�P,�EP�EPQ�J�у�]� U���}�H,�AV�u�R�Ѓ��    ^]�������������̡�}�P,�B����̡�}�P,�B����̡�}�P,�B����̡�}�P,�B ����̡�}�P,�B$����̡�}�P,�B(�����U���}�P,�R]�����������������U���}�P,�R��VW�E�P�ҋu����}�H�QV�ҡ�}�H$�QDV�ҡ�}�H$�QLVW�ҡ�}�H$�AH�U�R�Ћ�}�Q�J�E�P�у�_��^��]� �������U���}�H��D  ]��������������U���}�H��H  ]��������������U���}�H��L  ]��������������U���}�H�I]�����������������U���}�H�A]�����������������U���}�H�I]�����������������U���}�H�A]�����������������U���}�H�I]�����������������U���}�H���  ]��������������U���}�H�A]�����������������U���V�u�E�P���k�����}�Q$�J�E�P�у���u-��}�B$�PH�M�Q�ҡ�}�H�A�U�R�Ѓ�3�^��]Ë�}�Q�J�E�jP�у���u=�U�R��������u-��}�H$�AH�U�R�Ћ�}�Q�J�E�P�у�3�^��]Ë�}�B�HjV�у���u��}�B�HV�у����I�����}�Q$�JH�E�P�ы�}�B�P�M�Q�҃��   ^��]�����������U���}�H�A ]�����������������U���}�H�I(]�����������������U���}�H��  ]��������������U���}�H��   ]��������������U���}�H��  ]��������������U���}�H��  ]��������������U���}�H�A$��V�U�WR�Ћ�}�Q�u���BV�Ћ�}�Q$�BDV�Ћ�}�Q$�BLVW�Ћ�}�Q$�JH�E�P�ы�}�B�P�M�Q�҃�_��^��]������U���}�H���  ��V�U�WR�Ћ�}�Q�u���BV�Ћ�}�Q$�BDV�Ћ�}�Q$�BLVW�Ћ�}�Q$�JH�E�P�ы�}�B�P�M�Q�҃�_��^��]���U���}�H���  ]��������������U���<� ~SVW�E�    ��t�E�P�   �X������/��}�Q�J�E�P�   �ы�}�B$�PD�M�Q�҃��}��}�H�u�QV�ҡ�}�H$�QDV�ҡ�}�H$�QLVW�҃���t)��}�H$�AH�U�R����Ћ�}�Q�J�E�P�у���t&��}�B$�PH�M�Q�ҡ�}�H�A�U�R�Ѓ�_��^[��]���U���}�H�U���  ��VWR�E�P�ы�}�u���B�HV�ы�}�B$�HDV�ы�}�B$�HLVW�ы�}�B$�PH�M�Q�ҡ�}�H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡�}�H���   ��U���}�H���   V�uV�҃��    ^]�������������U���}�P�]���}�P�B����̡�}�P���   ��U���}�P�R`]�����������������U���}�P�Rd]�����������������U���}�P�Rh]�����������������U���}�P�Rl]�����������������U���}�P�Rp]�����������������U���}�P�Rt]�����������������U���}�P���   ]��������������U���}�P�Rx]�����������������U���}�P���   ]��������������U���}�P�R|]�����������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P�EPQ��  �у�]� �U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U��E��t ��}�R P�B$Q�Ѓ���t	�   ]� 3�]� U���}�P �E�RLQ�MPQ�҃�]� U��E��u]� ��}�R P�B(Q�Ѓ��   ]� ������U���}�P�R]�����������������U���}�P�R]�����������������U���}�P�R]�����������������U���}�P�R]�����������������U���}�P�R]�����������������U���}�P�R]�����������������U���}�P�E�R\P�EP��]� ����U���}�E�P�B ���$��]� ���U���}�E�P�B$Q�$��]� �����U���}�E�P�B(���$��]� ���U���}�P�R,]�����������������U���}�P�R0]�����������������U���}�P�R4]�����������������U���}�P�R8]�����������������U���}�P�R<]�����������������U���}�P�R@]�����������������U���}�P�RD]�����������������U���}�P�RH]�����������������U���}�P�RL]�����������������U���}�P�RP]�����������������U���}�P���   ]��������������U���}�P�RT]�����������������U���}�P�EPQ��  �у�]� �U���}�P���   ]��������������U���}�P���   ]��������������U���}�P�RX]����������������̡�}�P���   ��U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]��������������U���}�P���   ]�������������̡�}�P���   ��U���}�P���   ]�������������̡�}�P���   ���}�P���   ���}�P���   ��U���}�H���   ]��������������U���}�H��   ]��������������U���}�H�U�E��VWRP���  �U�R�Ћ�}�Q�u���BV�Ћ�}�Q�BVW�Ћ�}�Q�J�E�P�у�_��^��]������������U���}�H���  ]��������������U���}�P(�} �R8����P��]� �U���}�P�BdS�]VW��j ���Ћ�}�Q�����   h8�Fhc  V�Ћ�}���E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ�}�Q(�BHV���Ѕ�t ��}�Q(�E�R VP���҅�t�   �3��EP�R   ��_��^[]� ������U���V�E���MP�{���P���#�����}�Q�J���E�P�у���^��]� ���U��V�u���t��}�QP��Ѓ��    ^]���������̡�}�H��@  hﾭ���Y����������U��E��t��}�QP��@  �Ѓ�]����������������U���}�H���  ]��������������U���}�H��  ]�������������̡�}�H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�] ������u_^]Ã} tWj V��A ��_������F��}   ^]���U���}�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�\ ������u_^]�Wj V�VA ��_������F��}   ^]�������������U���}�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�\ ������u_^]�Wj V��@ ��_������F��}   ^]�������������U���}�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�[ ������u_^]�Wj V�V@ ��_������F��}   ^]�������������U���}�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�[ ������u_^]�Wj V��? ��_������F��}   ^]�������������U��M��t-�=�} t�y���A�uP��H ��]á�}�P�Q�Ѓ�]��������U��M��t-�=�} t�y���A�uP�H ��]á�}�P�Q�Ѓ�]��������U���}�H�U�R�Ѓ�]���������U���}�H�U�R�Ѓ�]���������U���}�E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��Y ������u_^]�Wj V�> ��_������F��}   ^]���������U���}�E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   ��}��t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��X ������u_^]�Wj V�= ��_������F��}   ^]����������U��E��w�   ��}��t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�@X ������u_^]�Wj V�= ��_������F��}   ^]�������U���}�H�U�R�Ѓ�]���������U���}�H�U�R�Ѓ�]���������U���}�H�U�R�Ѓ�]���������U���}�H�U�R�Ѓ�]���������U���}�Hp�]���}�Hp�h   �҃�������������U��V�u���t��}�QpP�B�Ѓ��    ^]���������U���}�Pp�EP�EPQ�J�у�]� U���}�Pp�EP�EPQ�J�у�]� U���}�Pp�EP�EPQ�J�у�]� U���}�Pp�EPQ�J�у�]� ���̡�}�HL���   ��U���}�H@�AV�u�R�Ѓ��    ^]�������������̡�}�HL�������U���}�H@�AV�u�R�Ѓ��    ^]�������������̡�}�PL���   Q�Ѓ�������������U���}�PL�EP�EPQ���   �у�]� �������������U���}V��HL���   V�҃���u��}�U�HL���   j RV�Ѓ�^]� ��}���   �ȋBP�Ћ�}���   �MP�BH��^]� �����̡�}�PL��(  Q�Ѓ�������������U���}�PL�EP�EPQ��,  �у�]� ������������̡�}�HL�Q�����U���}�H@�AV�u�R�Ѓ��    ^]��������������U���}�PL�E�R��VPQ�M�Q�ҋu��P���5r���M��Mr����^��]� ����U���}�PL�EPQ���   �у�]� �U���}�PL�EP�EPQ�J�у�]� ��}�PL�BQ�Ѓ���������������̡�}�PL�BQ�Ѓ���������������̡�}�PL�BQ�Ѓ����������������U���}�PL�EP�EP�EPQ�J �у�]� ������������U���}�PL�EPQ��4  �у�]� �U���}�PL�EP�EP�EPQ�J$�у�]� ������������U���}�PL�EP�EP�EP�EPQ�J(�у�]� �������̡�}�PL�B,Q�Ѓ���������������̡�}�PL�B0Q�Ѓ����������������U���}�PL�EP�EPQ��  �у�]� ������������̡�}�PL���   Q�Ѓ�������������U���}�PL�E��  ��VPQ�M�Q�ҋu��P���p���M��*p����^��]� ̡�}�PL�B4Q�Ѓ���������������̡�}�PL�B8j Q�Ѓ��������������U���}�PL���   ]��������������U���}�PL���   ]��������������U���}�PL���   ]��������������U���}�PL���   ]��������������U���}�PL���   ]��������������U���}�PL���   ]��������������U���}�PL���   ]��������������U���}�PL���   ]��������������U���}�PL���   ]��������������U���}�PL�EPQ�J<�у�]� ���̡�}�PL�BQ��Y�U���}�PL�EP�EPQ�J@�у�]� U���}�PL�Ej PQ�JD�у�]� ��U���}�PL�Ej PQ�JH�у�]� ��U���}�PL�EjPQ�JD�у�]� ��U���}�PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��tD  W�M�Q�U�R���dK  ���M�����6  ��t��}���   ��U�R�Ѓ�_^3�[��]Ë�}���   �J8�E�P�ы�}�����   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  �C  j�M�Q�U�R����J  �M��%6  ��}���   ��U�R�Ѓ�^��]�����������U���$��}�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��:C  j�E�P�M�Q���IJ  �M��5  ��}���   ��M�Q�҃�_^��]� ��U���$��}�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��B  j�E�P�M�Q����I  �M��!5  ��}���   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��TB  W�M�Q�U�R���DI  ���M����4  ��t+�u���i�����}���   ��U�R�Ѓ�_��^[��]� ��}���   �JL�E�P�ыu��P���������}���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��A  W�M�Q�U�R���H  ���M�����3  ��t+�u��������}���   ��U�R�Ѓ�_��^[��]� ��}���   �JL�E�P�ыu��P��������}���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}���@  W�M�Q�U�R����G  ���M����73  _^��[t��}���   ��U�R�������]Ë�}���   �J<�E�P���]���}���   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��$@  W�M�Q�U�R���G  ���M����2  ��t��}���   ��U�R�Ѓ�_^3�[��]Ë�}���   �J8�E�P�ы�}�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��t?  W�M�Q�U�R���dF  ���M�����1  ��t-��u��}����   ���^�U�R�Ѓ�_��^[��]� ��}���   �JP�E�P�ы�u�H��P�@�N��}�V���   �
�F�E�P�у�_��^[��]� �����̡�}�PL���   Q��Y��������������U���}�PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���}�PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}���=  W�M�Q�U�R����D  ���M����G0  ��t-��u��}����   ���^�U�R�Ѓ�_��^[��]� ��}���   �JP�E�P�ы�u�H��P�@�N��}�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��=  W�M�Q�U�R���D  ���M����w/  ��t-��u��}����   ���^�U�R�Ѓ�_��^[��]� ��}���   �JP�E�P�ы�u�H��P�@�N��}�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��D<  W�M�Q�U�R���4C  ���M����.  ��t-��u��}����   ���^�U�R�Ѓ�_��^[��]� ��}���   �JP�E�P�ы�u�H��P�@�N��}�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��t;  W�M�Q�U�R���dB  ���M�����-  ��t��}���   ��U�R�Ѓ�_^3�[��]Ë�}���   �J8�E�P�ы�}�����   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  �:  j�M�Q�UR����A  �M�&-  ��}���   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��O:  j�U�R�E�P���^A  �M��,  ��}���   �
�E�P�у�^��]� ��������U���$��}�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���9  j�E�P�M�Q����@  �M��1,  ��}���   ��M�Q�҃�_^��]� ��U���$��}�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J9  j�E�P�M�Q���Y@  �M��+  ��}���   ��M�Q�҃�_^��]� ��U���$��}�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���8  j�E�P�M�Q����?  �M��1+  ��}���   ��M�Q�҃�_^��]� ��U���$��}�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J8  j�E�P�M�Q���Y?  �M��*  ��}���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���7  j�U�R�E�P����>  �M��F*  ��}���   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}��t7  W�M�Q�U�R���d>  ���M�����)  ��t-��u��}����   ���^�U�R�Ѓ�_��^[��]� ��}���   �JP�E�P�ы�u�H��P�@�N��}�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��6  W�M�Q�U�R���=  ���M����)  ��t��}���   ��U�R�Ѓ�_^3�[��]Ë�}���   �J8�E�P�ы�}�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}���5  W�M�Q�U�R����<  ���M����W(  ��t��}���   ��U�R�Ѓ�_^3�[��]Ë�}���   �J8�E�P�ы�}�����   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U���$��}�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
5  j�E�P�M�Q���<  �M��q'  ��}���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��4  j�U�R�E�P���;  �M��'  ��}���   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��/4  j�U�R�E�P���>;  �M��&  ��}���   �
�E�P�у�^��]� ��������U���}�H���   ]��������������U���}�H���   ]�������������̡�}�H���   ���}�H���   ��U���}�H���   V�u�R�Ѓ��    ^]�����������U���}�H���   ]��������������U���}�HL�QV�ҋ���u^]á�}�H�U�ER�UP���  RV�Ѓ���u��}�Q@�BV�Ѓ�3���^]����������U���}�H�U�E���  R�U�� P�ERP�у�]������U���}�H���   ]��������������U���}�H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡�}�PL�BLQ�Ѓ���������������̡�}�PL�BPQ�Ѓ����������������U���}�PL�EP�EPQ�JT�у�]� U���}�PL�EPQ��  �у�]� �U���}�PL�EPQ���   �у�]� ̡�}�PL�BXQ�Ѓ����������������U���}�PL�EP�EP�EPQ�J\�у�]� ������������U���4��}SV��HL�QW�ҋ�3ۉ}�;��x  �M��!Z����}�E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ�}���   �BSSW���Ѕ���   ��}�QL�BW�Ћ���;���   ��    ��}���   �B(���ЍM�Qh�   ���u���  ������   �M�;���   ��}���   ���   S��;�tm��}���   �ȋB<V�Ћ�}���   ���   �E�P�у�;�t��}�B@�HV�у���;��\����}��M���   �M��YY����_^[��]� �}���}�B@�HW�ы�}���   ���   �M�Q�҃��M��y   �M��Y��_^3�[��]� �����̡�}�PL�B`Q�Ѓ���������������̡�}�PL�BdQ�Ѓ����������������U���}�PL�EPQ�Jh�у�]� ���̡�}�PL��D  Q�Ѓ������������̡�}�PL�BlQ�Ѓ����������������U���}�PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�EhphPh0h R�Q�U R�UR�UR�U���A�$�5�}�vLRP���   Q�Ѓ�4^]�  ������̡�}�PL���   Q�Ѓ�������������U���}�PL�EP�EP�EPQ��   �у�]� ���������U���}�PL��H  ]�������������̡�}�PL��L  ��U���}�PL��P  ]��������������U���}�PL��T  ]��������������U���}�PL�EP�EP�EP�EP�EPQ���   �у�]� �U���}�PL�EP�EP�EPQ���   �у�]� ���������U���}�PL�EP�EP�EP�EPQ��   �у�]� �����U���}�HL���   ]��������������U���}�HL���   ]��������������U���}�HL���   ]�������������̡�}�HL��  ���}�HL��@  ��h~Ph^� ��  ���������������U��Vh~j\h^� ����  ����t�@\��t
�MQV�Ѓ�^]� ������������U��� ��}V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\��}�QLjP���   ���ЋM��U�Rh=���M�}���  ����}���   ���   �U�R�Ѓ��M��u��  ��_^��]Ë�}���   ���   �E�P�у��M��u���  _�   ^��]����U��� ��}V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\��}�QLjP���   ���ЋM��U�Rh<���M�}��  ����}���   ���   �U�R�Ѓ��M��u��<  ��_^��]Ë�}���   ���   �E�P�у��M��u��  _�   ^��]����U���}�P8�EPQ�JD�у�]� ���̡�}�H8�Q<�����U���}�H8�A@V�u�R�Ѓ��    ^]�������������̡�}�H8�������U���}�H8�AV�u�R�Ѓ��    ^]��������������U���}�P8�EP�EP�EPQ�J�у�]� ������������U���}�P8�EP�EPQ�J�у�]� ��}�P8�BQ�Ѓ����������������U���}�P8�EPQ�J �у�]� ����U���}�P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U���}�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U���}�P8�EP�EPQ�J(�у�]� U���}�P8�EP�EP�EPQ�J,�у�]� ������������U���}�P8�EP�EP�EPQ�J�у�]� ������������U���}�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U���}�P8�EP�EPQ�J0�у�]� U���}�P8�EP�EP�EPQ�J4�у�]� ������������U���}�P8�EPQ�J8�у�]� ����U���}�H��x  ]��������������U���}�H��|  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H�A,]�����������������U���}�H�QV�uV�ҡ�}�H�Q8V�҃���^]�����̡�}�H�Q<�����U���}�H�I@]����������������̡�}�H�QD����̡�}�H�QH�����U���}�H�AL]�����������������U���}�H�IP]�����������������U���}�H��<  ]��������������U���}�H��,  ]��������������U���}�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡�}�H���   ���}�H���  ��U���}�H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U���}�H�A]�����������������U���}�H��\  ]��������������U���}�H�AT]�����������������U���}�H�AX]�����������������U���}�H�A\]����������������̡�}�H�Q`����̡�}�H�Qd����̡�}�H�Qh�����U���}�H�Al]�����������������U���}�H�Ap]�����������������U���}�H�At]�����������������U���}�H��D  ]��������������U���}�H��  ]��������������U���}�H�Ix]�����������������U���}�H��@  ]��������������U��V�u���²����}�H�U�A|VR�Ѓ���^]���������U���}�H���   ]��������������U���}�H��h  ]��������������U���}�H��d  ]��������������U���}�H���  ]�������������̡�}�H���   ��U���}�H��l  ]��������������U���}�H��   ]��������������U���}�H��  ]��������������U��V�u���RK����}�H���   V�҃���^]���������̡�}�H��`  ��U���}�H��  ]��������������U���}�H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U���}�H���  ]��������������U��U�E��}�H�E���   R���\$�E�$P�у�]�U���}�H���   ]��������������U���}�H���   ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���   ]��������������U���}�H���   ]��������������U���}�H���   ]��������������U���}�H���   ]��������������U���}�H���   ]��������������U���}�H���   ]��������������U���}�P���E�P�E�P�E�PQ���   �у����#E���]����������������U���}�P���E�P�E�P�E�PQ���   �у����#E���]����������������U���}�P���E�P�E�P�E�PQ���   �у����#E���]����������������U���}�H��8  ]��������������U��V�u(V�u$�E�@��}�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@��}�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U���}�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U���}�P0�EP�EP�EP�EPQ���   �у�]� ����̡�}�P0���   Q�Ѓ�������������U���}�P0�EP�EPQ���   �у�]� �������������U���}�P0�EP�EP�EP�EPQ���   �у�]� ����̡�}�P0���   Q�Ѓ������������̡�}�H0���   ��U���}�H0���   V�u�R�Ѓ��    ^]�����������U���}�H��H  ]��������������U���}�H��T  ]�������������̡�}�H��p  ���}�H���  ��U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H�U�E��X  ��VR�UPR�E�P�ыu�    �F    ��}���   �Qj PV�ҡ�}���   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M���D��P�E�hicMCP�k������M���D����}���   �JT�E�P�у���u(�u���jD����}���   ��M�Q�҃���^��]á�}���   �AT�U�R�Ћu��P���jD����}���   �
�E�P�у���^��]�������������U���}�H��  ]��������������U���}�H��\  ]��������������U���}�H�U��t  ��V�uVR�E�P�у���蓫���M��˪����^��]�����U���}�H�U���  ��VWR�E�P�ы�}�u���B�HV�ы�}�B�HVW�ы�}�B�P�M�Q�҃�_��^��]����������������U���}�H�U���  ��VWR�E�P�ы�}�u���B�HV�ы�}�B�HVW�ы�}�B�P�M�Q�҃�_��^��]����������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H�U�E��VWj R�UP�ERP��t  �U�R�Ћ�}�Q�u���BV�Ћ�}�Q�BVW�Ћ�}�Q�J�E�P�у�(_��^��]��U���}�H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    ��}���   j P�BV�Ћ�}���   �
�E�P�у�$��^��]���U���}�H��8  ]��������������U���  �Pg3ŉE��M�EPQ������h   R�`� ����|	=�  |#���}�H��0  hx�hF  �҃��E� ��}�H��4  ������Rh���ЋM�3̓��v ��]�������U���}�H��  ��V�U�WR�Ћ�}�Q�u���BV�Ћ�}�Q�BVW�Ћ�}�Q�J�E�P�у�_��^��]����U���}�H��  ��V�U�WR�Ћ�}�Q�u���BV�Ћ�}�Q�BVW�Ћ�}�Q�J�E�P�у�_��^��]����U���}�H��p  ��$�҅�trh���M��?����}�P�E�R4Ph���M��ҡ�}�P�E�R4Ph���M���j �E�P�M�hicMCQ������}���   ��M�Q�҃��M��?����]�U���}�H��p  ��$V�҅�u��}�H�u�QV�҃���^��]�Wh!���M���>����}�P�E�R4Ph!���M���j �E�P�M�hicMCQ������}���   �QHP�ҋu����}�H�QV�ҡ�}�H�QVW�ҡ�}���   ��U�R�Ѓ�$�M��>��_��^��]������U���}�H��p  ��$V�҅�u��}�H�u�QV�҃���^��]�Wh����M��,>����}�P�E�R4Ph����M���j �E�P�M�hicMCQ������}���   �QHP�ҋu����}�H�QV�ҡ�}�H�QVW�ҡ�}���   ��U�R�Ѓ�$�M���=��_��^��]������U���}�H��p  ��$�҅�u��]�Vh#���M��t=����}�P�E�R4Ph#���M���j �E�P�M�hicMCQ�������}���   �Q8P�ҋ��}���   ��U�R�Ѓ��M��U=����^��]���������������U���}�H��p  ��$�҅�u��]�Vhs���M���<����}�P�E�R4Phs���M���j �E�P�M�hicMCQ�W�����}���   �Q8P�ҋ��}���   ��U�R�Ѓ��M��<����^��]���������������U���}�H���  ]��������������U���}�H��@  ]��������������U���}�H���  ]��������������U��V�u���t��}�QP��D  �Ѓ��    ^]������U���}�H��H  ]��������������U���}�H��L  ]��������������U���}�H��P  ]��������������U���}�H��T  ]��������������U���}�H��X  ]��������������U���}�H��\  ]�������������̡�}�H��d  ��U���}�H��h  ]��������������U���}�H��l  ]�������������̡�}�H���  ��U���}�H�U���  ��VR�E�P�ыu��P���:���M��:����^��]�����U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H���  ]��������������U���}�H��$  ]��������������U���}�H��(  ]��������������U���}�H��,  ]�������������̡�}�H��0  ���}�H��<  ��U���}�H���  ]�������������̡�}�H���  ��U���}�H���  ]������������������������������U���}�H��  ]�������������̡�}�H��P  ���}���   ���   ��Q��Y��������U���}�H�A�U��� R�Ћ�}�Q�Jj j��E�h��P�ыUR�E�P�M�Q�[����}�B�P�M�Q�ҡ�}�H�A�U�R�Ћ�}�Q�J�E�P�у�,��]��h�}PhD �pz  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h�}jhD �y  ����t
�@��t]��3�]��������Vh�}j\hD ���ly  ����t�@\��tV�Ѓ���^�����Vh�}j`hD ���<y  ����t�@`��tV�Ѓ�^�������U��Vh�}jdhD ���	y  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�}jhhD ����x  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh�}jlhD ���x  ����t�@l��tV�Ѓ�^�������U��Vh�}h�   hD ���Vx  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�}h�   hD ���x  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�}jphD ���w  ����t�@p��t�MQV�Ѓ�^]� ��}^]� ��U��Vh�}jxhD ���yw  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�}jxhD ���9w  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�}jxhD ����v  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� ������������̋���������������h�}jhD �v  ����t	�@��t��3��������������U��V�u�> t+h�}jhD �cv  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h�}jhD �!v  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�}jhD ����u  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�}jhD ���u  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�}j hD ���\u  ����t�@ ��tV�Ѓ�^�3�^���Vh�}j$hD ���,u  ����t�@$��tV�Ѓ�^�3�^���U��Vh�}j(hD ����t  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�}j,hD ���t  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�}j(hD ���it  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�}j4hD ���t  ����t�@4��tV�Ѓ�^�3�^���U��Vh�}j8hD ����s  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�}j<hD ���s  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh�}jDhD ���\s  ����t�@D��tV�Ѓ�^�3�^���U��Vh�}jHhD ���)s  ����t�M�PHQV�҃�^]� U��Vh�}jLhD ����r  ����u^]� �M�PLQV�҃�^]� �����������U��Vh�}jPhD ���r  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�}jThD ���|r  ����u^Ë@TV�Ѓ�^���������U��Vh�}jXhD ���Ir  ����t�M�PXQV�҃�^]� U��Vh�}h�   hD ���r  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�}h�   hD ����q  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�}h�   hD ���vq  ����u^]� �M���   QV�҃�^]� �����U��Vh�}h�   hD ���6q  ����u^]� �M���   QV�҃�^]� �����U��Vh�}h�   hD ����p  ����u^]� �M���   QV�҃�^]� �����U��Vh�}h�   hD ���p  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh�}h�   hD �up  ����u��}�H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ�}�Q�u���BV�Ћ�}�Q�BVW�Ћ�}�Q�J�E�P�у�_��^��]��U��Vh�}h�   hD ����o  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�}h�   hD ���o  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�}h�   hD ���Vo  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�}h�   hD ���o  ����t���   ��t�MQ����^]� 3�^]� �Vh�}h�   hD ����n  ����t���   ��t��^��3�^����������������U��Vh�}h�   hD ���n  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�}h�   hD ���Fn  ����t���   ��t�MQ����^]� ��������U��Vh�}h�   hD ���n  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh�}h�   hD ���m  ����t���   ��t��^��3�^����������������VW��3����$    �h�}jphD �om  ����t�@p��t	VW�Ѓ����}�8 tF��_��^�������U��SW��3�V��    h�}jphD �m  ����t�@p��t	WS�Ѓ����}�8 tqh�}jphD ��l  ����t�@p��t�MWQ�Ѓ������}h�}jphD �l  ����t�@p��t	WS�Ѓ����}V���7�����tG�]����E^��t�8��~=h�}jphD �nl  ����t�@p��t	WS�Ѓ����}�8 u_�   []� _3�[]� ����������U��Vh�}j\hD ���l  ����t3�@\��t,V��h�}jxhD ��k  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�}j\hD ���k  ����t3�@\��t,V��h�}jdhD �k  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�}j\hD ���Vk  ����tG�@\��t@V�ЋEh�}jdhD �E��E�    �E�    � k  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�}j\hD ����j  ����t\�@\��tUV��h�}jdhD �j  ����t�@d��t
�MQV�Ѓ�h�}jhhD �j  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�}j\hD ���Ij  ������   �@\��t~V��h�}jdhD �#j  ����t�@d��t
�MQV�Ѓ�h�}jhhD ��i  ����t�@h��t
�URV�Ѓ�h�}jhhD ��i  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh�}jthD ���i  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�}j`hD �^i  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh�}���_�����^��]� ������U���Vh�}h�   hD ���i  ����tR���   ��tH�MQ�U�R���ЋuP������h�}j`hD ��h  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t��}���   P�B@��]� �E��t��}���   P�BD��]� ��}���   R�PD��]� �����U���}�P@�Rd]�����������������U���}�P@�Rh]�����������������U���}�P@�Rl]�����������������U���}�P@�Rp]�����������������U���}���   ���   ]�����������U���}���   ���   ]����������̡�}�P@�Bt����̡�}�P@�Bx�����U���}�P@�R|]����������������̡�}�P@���   ���}���   �Bt��U���}�P@���   ]�������������̡�}�P@���   ��U���}�P@���   ]��������������U���}�P@���   ]��������������U���}�P@���   ]��������������U���}�P@���   ]��������������U���}V��H@�QV�ҋM����t��#�����}�Q@P�BV�Ѓ�^]� �̡�}�PH���   Q�Ѓ�������������U���}�P@�EPQ�JL�у�]� ���̡�}�P@�BHQ�Ѓ����������������U���}�P@�EP�EP�EPQ�J�у�]� ������������U���}�P@�EPQ�J�у�]� ����U���}�P@�EP�EPQ�J�у�]� U���}�P@�EPQ�J �у�]� ����U���}���   �R]��������������U���}���   �R]��������������U���}���   �R ]��������������U���}���   ���   ]�����������U���}���   ��D  ]�����������U���}�E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U���}���   ���   ]����������̡�}���   �B$���}�H@�Q0�����U���}�H@�A4j�URj �Ѓ�]����U���}�H@�A4j�URh   @�Ѓ�]�U���}�H@�U�E�I4RPj �у�]�̡�}�H|�������U��V�u���t��}�Q|P�B�Ѓ��    ^]��������̡�}�H|�Q �����U��V�u���t��}�Q|P�B(�Ѓ��    ^]��������̡�}�H@�Q0�����U��V�u���t��}�Q@P�B�Ѓ��    ^]���������U���}�H@���   ]��������������U��V�u���t��}�Q@P�B�Ѓ��    ^]��������̡�}�PH���   Q�Ѓ�������������U���}�PH�EPQ��d  �у�]� �U���}�H �IH]�����������������U��}qF uHV�u��t?��}���   �BDW�}W���Ћ�}�Q@�B,W�Ћ�}�Q�M�Rp��VQ����_^]����������̡�}�P@�BT�����U���}�P@�RX]�����������������U���}�P@�R\]����������������̡�}�P@�B`�����U���}�H��T  ]��������������U���}�H@�U�A,SVWR�Ћ�}�Q@�J,���EP�ы�}�Z��h��hE  �΋��v��Ph��hE  ���d��P��T  �Ѓ�_^[]����U���}�PT�EP�EPQ�J�у�]� U���}�PT�EPQ�J�у�]� ����U���}�PT�EPQ�J�у�]� ����U���}�PT�E�R<��PQ�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U���}�HT�]��U���}�H@�AV�u�R�Ѓ��    ^]�������������̡�}�HT�hG  �҃�������������U���}�H@�AV�u�R�Ѓ��    ^]�������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�BQ�Ѓ����������������U���}�PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U���}�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U���}�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U���}�PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U���}�PX�EPQ�J�у�]� ����U���}�PX�EPQ�J�у�]� ����U���}�PX�EPQ�J�у�]� ����U���}�PX�EPQ�J�у�]� ����U���}�PX�EPQ�J$�у�]� ����U���}�PX�EPQ�J �у�]� ����U���}�PD�EP�EPQ�J�у�]� U���}�HD�U�j R�Ѓ�]�������U���}�H@�AV�u�R�Ѓ��    ^]��������������U���}�HD�	]��U���}�H@�AV�u�R�Ѓ��    ^]��������������U���}�HD�U�j R�Ѓ�]�������U���}�H@�AV�u�R�Ѓ��    ^]��������������U���}�U�HD�Rh'  �Ѓ�]����U���}�H@�AV�u�R�Ѓ��    ^]�������������̡�}�HD�j h�  �҃�����������U���}�H@�AV�u�R�Ѓ��    ^]�������������̡�}�HD�j h:  �҃�����������U���}�H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E���}���   �R�E�Pj�����#E���]�̡�}�HD�j h�F �҃�����������U���}�H@�AV�u�R�Ѓ��    ^]�������������̡�}�HD�j h�_ �҃�����������U���}�H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E���}�E�    ���   �R�E�Pj������؋�]� ̡�}�PD�B$Q�Ѓ���������������̡�}�PD�B(Q�Ѓ���������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�B(Q�Ѓ���������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�B(Q�Ѓ���������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�B(Q�Ѓ���������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�B(Q�Ѓ���������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�B(Q�Ѓ���������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�B(Q�Ѓ���������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�B(Q�Ѓ���������������̡�}�PD�BQ�Ѓ���������������̡�}�PD�B(Q�Ѓ���������������̡�}�PD�BQ�Ѓ����������������U���}�H �Ah]�����������������U���}�H@�AV�u�R�Ѓ��    ^]�������������̡�}�H �������U��V�u���t��}�Q P�B�Ѓ��    ^]���������U���}�P �EPQ�J4�у�]� ����U���}�P �EPQ�J�у�]� ����U���}�P �EPQ�J�у�]� ���̡�}�P �BQ��Y�U��V�uW����������}�H �QVW�҃�_��^]� �����U���}�P �EPQ�J �у�]� ���̡�}�P �B,Q�Ѓ���������������̡�}�P �B0Q�Ѓ���������������̡�}�H\�������U���}�H\�AV�u�R�Ѓ��    ^]�������������̡�}�P\�BQ�Ѓ���������������̡�}�P\�BQ�Ѓ����������������U���}�P\�EPQ�J�у�]� ����U���}�P\�EP�EPQ�J�у�]� U���}�P\�EPQ�J�у�]� ���̡�}�P\�BQ�Ѓ����������������U���}�P\�EPQ�J �у�]� ����U���}�P\�EP�EPQ�J$�у�]� U���}�P\�EP�EP�EPQ�J(�у�]� ������������U���}�P\�EPQ�J0�у�]� ����U���}�P\�EPQ�J@�у�]� ����U���}�P\�EPQ�JD�у�]� ����U���}�P\�EPQ�JH�у�]� ���̡�}�P\�B4Q�Ѓ����������������U���}�P\�EP�EPQ�J8�у�]� U���}�P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu��������}�H\�QV�҃���S���ۏ��3���~=��I ��}�H\�U�R�U��EP�A(VR�ЋM��Q��訏���U�R��蝏��F;�|�_^[��]� ���������������U���VW�}�E��P�������}� ��   ��}�Q\�BV�Ѓ��M�Q��������E���t]S3ۅ�~H�I �UR��襋���E�P��蚋���E;E�!����}�Q\P�BV�ЋE@��;E��E~�C;]�|�[_�   ^��]� _�   ^��]� U���}�E�PH�B���$Q�Ѓ�]� ���������������U���}�PH�EPQ���   �у�]� �U���}�PH�EPQ���  �у�]� �U���}�PH�EPQ���  �у�]� �U���}�PH�EP�EPQ��  �у�]� �������������U���}�PH�EP�EPQ��  �у�]� ������������̡�}�PH���  Q�Ѓ�������������U���}�PH�EPQ���  �у�]� ̡�}�PH���   j Q�Ѓ�����������U���}�PH�EPj Q���   �у�]� ��������������̡�}�PH���   jQ�Ѓ�����������U���}�PH�EPjQ���   �у�]� ��������������̡�}�PH���   jQ�Ѓ����������U���}�PH�EPjQ���   �у�]� ���������������U���}�PH�EP�EPQ���   �у�]� �������������U���}�PH�EP�EPQ���   �у�]� ������������̡�}�PH���   Q�Ѓ�������������U���}�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP�������������t�E��}�QH���   PVW�у���_^]� �����U��EVW���MPQ�����������t�M��}�BH���   QVW�҃���_^]� ̡�}�PH���   Q�Ѓ������������̡�}�PH���   Q�Ѓ�������������U���}�PH�EPQ���   �у�]� �U���}�PH�EPQ���   �у�]� �U���}�PH�EP�EPQ��8  �у�]� �������������U���}�PH�EP�EPQ��   �у�]� ������������̡�}�PH���  Q�Ѓ������������̡�}�PH���  Q�Ѓ������������̡�}�PH���  Q�Ѓ������������̡�}�PH��  Q�Ѓ������������̡�}�PH��  Q�Ѓ�������������U���}�PH�EP�EPQ��  �у�]� �������������U���}�PH�EP�EP�EPQ��   �у�]� ���������U���}�PH�EP�EP�EP�EPQ��|  �у�]� �����U���}�PH�EPQ��  �у�]� ̡�}�PH��T  Q�Ѓ�������������U���}�PH�EP�EPQ��  �у�]� �������������U���}�PH�EPQ��8  �у�]� �U���}�PH�EPQ��<  �у�]� �U���}�PH�EPQ��@  �у�]� �U���}�PH�EP�EP�EPQ��D  �у�]� ��������̡�}�PH��L  Q��Y��������������U���}�PH�EPQ��H  �у�]� ̡�}V��H@�Q,WV�ҋ�}�Q��j �ȋ��   h�  �Ћ�}�QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡�}�P@�B,Q�Ћ�}�Q��j �ȋ��   h�  �������U���}�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U���}�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U���}�PH�EP�EP�EPQ��   �у�]� ��������̡�}�HH��  ��U���}�HH��  ]��������������U���}�E�PH��$  ���$Q�Ѓ�]� �����������̡�}�PH��(  Q�Ѓ�������������U���}�PH�EP�EPQ��,  �у�]� �������������U���}�E�PH�EP�E���$PQ��0  �у�]� ���̡�}�PH���  Q�Ѓ������������̡�}�PH��4  Q�Ѓ������������̋��     �������̡�}�PH���|  jP�у���������U���}�UV��HH��x  R��3Ƀ������^��]� ��̡�}�PH���|  j P�у��������̡�}�PH��P  Q�Ѓ������������̡�}�PH��T  Q�Ѓ������������̡�}�PH��X  Q�Ѓ�������������U���}�PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡�}�PH��`  Q�Ѓ�������������U���}�PH�EPQ��d  �у�]� �U���}�E�PH��h  ���$Q�Ѓ�]� ������������U���}�E�PH��t  ���$Q�Ѓ�]� ������������U���}�E�PH��l  ���$Q�Ѓ�]� ������������U���}�PH�EPQ��p  �у�]� �U���}�PH�EP�EP�EP�EPQ���  �у�]� �����U���}�PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U���}�E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E��}�HH�E���   R�U���$P�ERP�у�]����������������U���E�M�����  �M;�|�M;�~��]�����������U���}�PH�E���   Q�MPQ�҃�]� ������������̡�}�PH���   Q��Y�������������̡�}�PH���   Q�Ѓ������������̡�}�PH���   Q��Y��������������U���}�PH�EP�EPQ���   �у�]� �������������U���}�PH�EP�EP�EP�EP�EPQ���  �у�]� ̡�}�PH��t  Q��Y�������������̋�� ���@    ������}�Pl�A�JP��Y��������U���}V��Hl�V�AR�ЋE����u
�   ^]� ��}�Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË�}�QlP�B�Ѓ�������U���}�Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E��}�HH�ER�U���$P���  R�Ѓ�]����U���}�HH���  ]��������������U���}�HH���  ]��������������U��U0�E(��}�HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U���}�HH���  ]��������������U���}�E�PH�EP���$Q���  �у�]� ��������U���SV��������؉]����   �} ��   ��}�HH��p  j h�  V�҃��E��u
^��[��]� �MW3��}����������   �]��I �E�P�M�Q�MW������ta�u�;u�Y�I ������u�E�������L�;Ht-��}�Bl�S�@����QR�ЋD������t	�M�P�s���F;u�~��}��MG�}��>���;��v����]�_^��[��]� ^3�[��]� ��������������U�����}SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u��}�HH���  �'��u��}�HH���  ���uš�}�HH���  S�ҋȃ��E��t�W������}�HH���   h�  S3��҃����  ���_�u����    ��}�Hl�U�B�IWP�ы�������   ��}�F�J\�UP�A,R�Ѓ���t�K�Q�M�%�����}�F�J\�UP�A,R�Ѓ���t�K�Q�M������E��;Pt&�F��}�Q\�J,P�EP�у���t	�MS�������}�v�B\�M�P,VQ�҃���t�M�CP������}�QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U���}�HH���   ]�������������̡�}�PH���   Q��Y��������������U���}�HH���  ]��������������U���}��P���   V�uW�}���$V�����E������At���E������z����؋�}�Q�B,���$V����_^]����������������U���0���}�U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١�}�]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U���}�HH�]��U���}�H@�AV�u�R�Ѓ��    ^]�������������̡�}�HH�h�  �҃�������������U���}�H@�AV�u�R�Ѓ��    ^]��������������U���}�HH�Vh  �ҋ�������   �EPh�  � �������t]��}�QHj P���   V�ЋMQh(  ���������t3��}�JH���   j PV�ҡ�}���   �B��j j���Ћ�^]á�}�H@�QV�҃�3�^]�������U���}�H@�AV�u�R�Ѓ��    ^]��������������U���}�HH�Vh�  �ҋ�����u^]á�}�HH�U�E��  RPV�у���u��}�B@�HV�у�3���^]�������U���}�H@�AV�u�R�Ѓ��    ^]��������������U���}�HH�I]�����������������U���}�H@�AV�u�R�Ѓ��    ^]��������������U���}�PH�EPQ���  �у�]� �U���}�PH�EPQ���  �у�]� ̡�}�PH���  Q�Ѓ�������������U���}�HH���  ]��������������U���}�E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡�}�PH���  Q�Ѓ�������������U���}�PH�EP�EPQ���  �у�]� ������������̡�}�PH��  Q�Ѓ�������������U���}�PH�EP�EP�EPQ���  �у�]� ��������̡�}�PH���  Q�Ѓ������������̡�}�PH���  Q�Ѓ�������������U���}�PH�EPQ��  �у�]� �U���}�PH�EPQ��  �у�]� ̋������������������������������̡�}�HH���  ��U���}�HH���  ]��������������U���}�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U���}�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡�}�PH��,  Q�Ѓ�������������U���}�PH�EPQ��X  �у�]� ̡�}�PH��\  Q�Ѓ�������������U���}�HH��0  ]��������������U���}��W���HH���   j h�  W�҃��} u�   _��]� Vh�  ������������   ��}�HH���   j VW�҃��M��s�����}�P�E�R0Ph�  �M����E��}�P�B,���$h�  �M��Ћ�}�Q@�J(j �E�PV�у��M��|���^�   _��]� ^3�_��]� �����U��S�]�; VW��u7��}�U�HH���   RW�Ѓ���u��}�QH���   jW�Ѓ���t�   �����   ��}�QH���   W�Ѓ��} u(��}�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;��}�U�HH�ER�USP���  VRW�Ћ�}���   �B(�����Ћ���uŃ; u��}�QH���   W�Ѓ���t3���   �W��u1��}�QH���   �Ћ�}�E�QH���   PW�у�_^[]� ��}�BH���   �у��} u0��}�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ��}�QH�h  �Ћ؃���u_^[]� ��}���   �u�Bx���Ћ�}���   P�B|���Ѕ�tU��}�E�QH�MP�Ej Q���  VPW�у���t��}���   �ȋBHS�Ћ�}���   �B(���Ћ���u�_^��[]� ��������������U��EV���u��}�HH���  �'��u��}�HH���  ���u��}�HH���  V�҃���u3�^]� P�EP���>���^]� ���������U���D��}�HH���   S�]VWh�  S�ҋ��}�HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��.
  ��}���   �B���Ћ�}=�  ��  �QH���   Wh:  S�Ћ�}�QH�E����   h�  S�Ћ�}�QHW�����   h�  S�uԉ}��Ћ�}�QH�E苂  S�Ћ�}�QH�EЋ��  S�Ѓ�(�E��E�����~~�M���M�I �MЅ�tMj�W��m  ���t@�@�Ẽ|� �4�~����%�������;�u/����v  ;E�~�E؋��v  E���E�;Pu�E���E��E�G;}�|��}� tv�u�j S���{�������  ���������tV�������}�;�uK��}�H���  �4�h����h�  V�҃��E���N  �M�PVP�}���P�w}  ����}ܡ�}�H���  �4�h����h�  V�҃��E����  �M�3�;�t;�tVQP��  ���E�;�~-��}�Qh����h�  P���   �Ѓ��E�;���  ��}�E��QH��  j�PS�у�����  �u�;�tjS���]������{  ��������E���}��}�BH���   Wh�  S�у�3�9}ԉE�}��`  �}���}Ȑ�MЅ��R  �U�j�R��k  ����>  �M̍@�|� ���]�~����%�������9E���  ���t  �E�3�3�9C�E܉M���   ��$    �����������tk�]��}������������ϋ9�<��}�@�҉��y�]��|��]�@@�z�<��y�]��|��]�@@�z�<��I�}��]�@���M��}�@����@�M�A;K�M��t����E؅��9  �+U�j��PR�M���X  �M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$�D��U����4�"�M����t��U����t�
�M����t�M���;]�|��E܃�F;]؉M��	����U�;U��
  �U�R��q���E�P�q���M�Q�q����_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���P�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@��;EԉE��}�������U�R�o���E�P�o�����  ���   �B����=  ��  ��}�QH���   j h(  S�Ћ�}�QH�����   h(  S�ЋЃ�3��U؅�~'����    �ǅ�t�|� t�4N��tN�@;�|�u��u܋�}�Q���  �4v�h����hK  V�Ѓ��E�����   �M��t��tVQP��  ���u؋�}�Q���  �h����hP  V�Ѓ��E���tP��t��tVWP�f�  ���M����+�}�RH��PQ�E���   S�Ѓ���u�M�Q�Rn���U�R�In����_^3�[��]á�}�HH���   j h�  S�҉E���}�HH���   j h(  S��3�3���3�9]؉E��}ĉ]��7  �U��څ��  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�F@F����;�|��}ă|� ts�U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�F�v�Ћ��A�B�A�B�A�B�A�B�I�J�U�F<ډ}�C;]؉]�������M�3�3�;�~�U����$    ��t���   @;�|��U�R�l�����E�P�{l����_^�   [��]Ï�������������������U��E� �M+]� ���������������U��V��V�����}�Hl�AR�Ѓ��Et	V�Do������^]� ����������h�}Ph�f �*  ���������������U���Vh�}h�   h�f ����)  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh�}h�   h�f ���V)  ����t���   ��t�M�UQ�MRQ����^]� U���Vh�}h�   h�f ���)  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh�}h�   h�f ���(  ����t���   ��t�M�UQ�MRQ����^]� U��Qh�}h�   h�f �H(  ����t���   �E���t�EP�U�����]��@���]�������������U���h�}h�   h�f ��'  3Ƀ�;�tK9��   tC�E���   ���M��$Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]ËE�   � �  �P�P�H�H�H��]��U��h�}h�   h�f �i'  ����t���   ��t]��]����U��h�}h�   h�f �9'  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h�}h�   h�f ��&  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h�}h�   h�f �y&  ����t���   ��t]��3�]��U���Vh�}h�   h�f �E&  ����tZ���   ��tP�M�UWQR�M�Q�Ћ�}�u���B�HV�ы�}�B�HVW�ы�}�B�P�M�Q�҃�_��^��]á�}�H�u�QV�҃���^��]����������h�}h�   h�f �%  ����t���   ��t��3��������U��h�}h�   h�f �y%  ����t���   ��t]��]����U��M��U+u&�A+Bu�A+Bu�A+Bu�A+Bu�A+B]����������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���h�}�   h�   h�f �E��  �E��E��E�    �E�    �E�    ��"  ����t���   ��t	�M�Q�Ѓ��UR�E�P��������]��U��E��u��}�MP�EPQ������]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h0�j;h ~j�=h������t
W���~F���3��F��u_^]� �~ t3�9_��^]� ��}�H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ��}�H<�Q��3Ʌ����^��������������̃y t�   ËA��uË�}�R<P��JP�у��������U����u��}�H�]� ��}�J<�URP�A�Ѓ�]� ���������������U���}��u��}�H�]Ë�}�J<�URP�A�Ѓ�]�U���}��$V��u��}�H�1���}�J<�URP�A�Ѓ�����}�Q�J�E�SP�ы�}�B�P�M�QV�ҡ�}�H�A�U�R�Ћ�}�Q�Jj j��E�ht�P�ы�}�B�@@�� j �M�Q�U�R�M��Ћ�}�Q�J���E�P���у���[t.��}�B�u�HV�ы�}�B�P�M�Q�҃���^��]á�}�P�E��RHjP�M��ҡ�}�P�E�M��RLj�j�PQ�M��ҡ�}�H�u�QV�ҡ�}�H�A�U�VR�Ћ�}�Q�J�E�P�у���^��]���������������U���}��$SV��u��}�H�1���}�J<�URP�A�Ѓ�����}�Q�J�E�P�ы�}�B�P�M�QV�ҡ�}�H�A�U�R�Ћ�}�Q�Jj j��E�ht�P�ы�}�B�@@�� j �M�Q�U�R�M��Ћ�}�Q�J���E�P���у���t/��}�B�u�HV�ы�}�B�P�M�Q�҃���^[��]á�}�P�E��RHjP�M��ҡ�}�P�E�M��RLj�j�PQ�M��ҡ�}�H�A�U�R�Ћ�}�Q�Jj j��E�ht�P�ы�}�B�@@��j �M�Q�U�R�M��Ћ�}�Q�J���E�P���у����3�����}�P�E��RHjP�M��ҡ�}�P�E�M��RLj�j�PQ�M��ҡ�}�H�u�QV�ҡ�}�H�A�U�VR�Ћ�}�Q�J�E�P�у���^[��]����������������U���}��$SV��u��}�H�1���}�J<�URP�A�Ѓ�����}�Q�J�E�P�ы�}�B�P�M�QV�ҡ�}�H�A�U�R�Ћ�}�Q�Jj j��E�ht�P�ы�}�B�@@�� j �M�Q�U�R�M��Ћ�}�Q�J���E�P���у���t/��}�B�u�HV�ы�}�B�P�M�Q�҃���^[��]á�}�P�E��RHjP�M��ҡ�}�P�E�M��RLj�j�PQ�M��ҡ�}�H�A�U�R�Ћ�}�Q�Jj j��E�ht�P�ы�}�B�@@��j �M�Q�U�R�M��Ћ�}�Q�J���E�P���у����3�����}�P�E��RHjP�M��ҡ�}�P�E�M��RLj�j�PQ�M��ҡ�}�H�A�U�R�Ћ�}�Q�Jj j��E�ht�P�ы�}�B�@@��j �M�Q�U�R�M��Ћ�}�Q�J���E�P���у����������}�P�E��RHjP�M��ҡ�}�P�E�M��RLj�j�PQ�M��ҋu�E�P���sv����}�Q�J�E�P�у���^[��]�������U���}��$SV��u��}�H�1���}�J<�URP�A�Ѓ�����}�Q�J�E�P�ы�}�B�P�M�QV�ҡ�}�H�A�U�R�Ћ�}�Q�Jj j��E�ht�P�ы�}�B�@@�� j �M�Q�U�R�M��Ћ�}�Q�J���E�P���у���t/��}�B�u�HV�ы�}�B�P�M�Q�҃���^[��]á�}�P�E��RHjP�M��ҡ�}�P�E�M��RLj�j�PQ�M��ҡ�}�H�A�U�R�Ћ�}�Q�Jj j��E�ht�P�ы�}�B�@@��j �M�Q�U�R�M��Ћ�}�Q�J���E�P���у����3�����}�P�E��RHjP�M��ҡ�}�P�E�M��RLj�j�PQ�M��ҡ�}�H�A�U�R�Ћ�}�Q�Jj j��E�ht�P�ы�}�B�@@��j �M�Q�U�R�M��Ћ�}�Q�J���E�P���у����������}�P�E��RHjP�M��ҡ�}�P�E�M��RLj�j�PQ�M���j ht��M��t����}�P�R@j �E�P�M�Q�M��҅���}�H�A�U�R���Ѓ���t/��}�Q�u�BV�Ћ�}�Q�J�E�P�у���^[��]Ë�}�M��B�PHjQ�M��ҡ�}�P�E�M��RLj�j�PQ�M��ҋu�E�P���;s����}�Q�J�E�P�у���^[��]���������������U���}�H<�A]����������������̡�}�H<�Q�����V��~ u>���t��}�Q<P�B�Ѓ��    W�~��t����;��W�\�����F    _^��������U���V�E�P���~M����P��������M���;����^��]��̃=�} uK��}��t��}�Q<P�B�Ѓ���}    ��}��tV���`;��V�
\������}    ^������������U���8��}�H�AS�U�V3�R�]��Ћ�}�Q�JSj��E�hx�P�ы�}�B<�P�M�Q�ҋ��}�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��h  �M�Q�U�R�M��  ����   W�}�}���   ��}���   �U��ATR�Ћ�����tB��}�Q�J�E�P���у��U�Rj�E�P���q����}�Q�ȋBxW���E���t�E� ��t��}�Q�J�E�P����у���t��}�B�P�M�Q����҃��}� u"�E�P�M�Q�M���  ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3ۉ]�;�u_��}�H�A�U�R�Ћ�}�Q�JSj��E�hx�P�ы�}�B<�P�M�Q�ҋ��}�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]���  �M�Q�U�R�M��1  ���p  W�}��I �E����   ��}���   �U��ATR�Ћ�������   ��}�Q�J�E�P���ы�}�B���   ���M�Qj�U�R���Ћ�}�Q�J���E�P�ы�}�B�P�M�QV�ҡ�}�H�A�U�R�Ћ�}�Q�Bx��W�M����E��t�E ��t��}�Q�J�E�P����у���t��}�B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*��}���   P�BH�Ћ�}�Q���ȋBxW�Ѕ�t"�M�Q�U�R�M���  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��3  �EP�M�Q�M�u��u�}  ����   �u���E���tA��t<��uZ��}���   �M�PHQ�ҋ�}�Q���ȋBxV�Ѕ�u-�   ^��]Ë�}���   �E�JTP��VP�[�������uӍUR�E�P�M���  ��u�3�^��]����������V��~ u>���t��}�Q<P�B�Ѓ��    W�~��t���6��W�TW�����F    _^�������̋�� ����������������������̅�t��j�����̡�}�P��  ���}�P��(  ��U���}�P��   ��V�E�P�ҋuP����5���M��6����^��]� ��������̡�}�P��$  ��U���}�H��  ]��������������U���}�H���  ]�������������̡�}�H��  ��U���}�H���  ]��������������U���}�H��x  ]��������������U���}�H��|  ]��������������U���EV�����t	V��U������^]� �������������̸   � �������̸   @� �������̸   � �������̸   � ��������U���}�H�QV�uV�҃���^]� �3�� �����������3�� �����������U����   h�   ��@���j P�Ԕ  �M�Eh�   ��@���R�M��MPQjǅ`���    �~���� ��]���U����   V�u��u3�^��]�h�   ��@���j P�u�  �M�U�Eh�   �M���@���Q�U��U��@����ERPj��`���ǅD���Т�E�'�E����E����E��'�E� ��E�p��E����}���� ^��]�������������U���   SV�u(3ۉ]���u��}�H�A�UR�Ѓ�^3�[��]Ë�}�Q�B<W�M3��Ѕ��'  ��Y  �E���tq�MQ�M��2��Wh���M��j��P�M��2���u�Wj��U�R�E�P��\���Q�_?�D����P��x���R�E6����P�E�P�86����P���[  �E���t�E� �� t�M�����2����t��x�������2����t��\�������2����t�M̃���z2����t��}�Q�J�E�P����у���t�M��P2���}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R�X  ����E$�M�UVP�Ej QRP�����������}�Q�J�EP�у���_^[��]���������������̋�`����������̋�`����������̋�`����������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V���W  �����   �ESP�M���/����}�Q�J�E�P�ы�}�B�Pj j��M�h��Q�҃��E�P�M��/��j j��M�Q�U�R��d���P��A����P�M�Q�w3����P�U�R�j3�����P�?X  ���M�����/���M���/����d�����/���M���/����}�H�A�U�R�Ѓ��M��/����[t	V�OV  ����^��]� ���U��EVP����_  �����^]� �����Q�V  Y���������U��E�M�U�H4�M�P �U��M�@Т�@8'�@<��@@���@Dp��@H ��@L���@P��@l '�@X�'�@\�&�@`p'�@d0'�@T�'�@h`'�@p�&�@t ��P0�H(�@,    ]��������������U���   h�   ��`���j P��  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�x����8��]��������������̋�` ����������̋�`@����������̋�`����������̋�`�����������U���EV���V��������Au��}�H��0  h��j,�����^��^]� �����U���W������G���U����������A�  ������A��   ���������AuR������AuKV�����  �����  �ȅ�u��^����__��]Ëƙ����ʅ�u�u��E�^������__��]���������Au������=����������Au6�����������U������G�����_��������Au�����U����_�
����������ݭ  �E����U������������A{���������__��]�������������__��]����U�����V�E��������At�����������Au��������������$蚥  ���������^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3������;���W���$���!�  ��E������$��  �V����������Au��}�H��0  h��j�����^����_u������������^]� ���U������EV�ы�������z!��}�؋H��0  h��j5�����U������$�y�  �]��F�$�k�  �}��$�`�  ��E�$�S�  �^�����&���^��]� ���������������U���}���   �BXQ�Ѓ���u]� ��}�Q|�M�RQ�MQP�҃�]� ���U���}���   �BXQ�Ѓ���u]� ��}�Q|�M�R8Q�MQP�҃�]� ���U��EV��j ���}�Qj j P�B�ЉF����^]� ��̡�}Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ��}�Q�MP�EP�Q�JP�у��F�   ^]� ����U��M��P]����U��M��P]����U��M��P]����V������F    ��}�HP�h��Vh��h���҉F����^����������̃y ���u��}�PP�A�JP��Y��U��A��u]� ��}�QP�M�Rj Q�MQP�҃�]� ��U��A��t��}�QP�M�RQP�҃�]� ������������U��A��t��}�QP�M�RQP�҃�]� �����������̡�}�HP���   ��U���}�HP���   ]�������������̡�}�HP�QP�����U���}�HP�AT]����������������̋��     �@    �V����t)��}�QPP�BL�Ћ�}�QP��J<P�у��    ^�������������U��SV�ً3�W;�t��}�QPP�B<�Ѓ��3�s�}�Eh��W�C��}�QP�J8h��h��P�EP�у�9u�~M�I ���z u!���@   ��}�QP���H�RQ�҃���}�HP��A@VR�Ћ�F��;u�A|�3�9_^��[]� ��������U��SVW��3�9w~<�]��}�HP��A@VR�Ѓ���t-��}�QPj SjP�B�Ѓ���tF;w|�_^�   []� ��}�QP��JLP�у�_^3�[]� �����������̡�}�PP��JDP�у�������������̡�}�PP��JHP��Y��������������̡�}�PP��JLP��Y���������������U��U�E�@R�URP�I���]� �����U��V��~ ���u��}�HP�V�AR�Ѓ��Et	V�F������^]� ����U��E��u�E�M�~�~�   ]� �����������U��EHV����   �$����   ^]á~@�~��uT�EP�7�����=�.  }�����^]Ëu��t�h�jmh ~j��F������t ���]$��� ~��tV���l(���   ^]�� ~    �   ^]ËM�UQR蕥���������H^]�^]�@����-~u.�b����M���� ~��t����$��V�E����� ~    �   ^]Ã��^]ÍI ��9�@�����U��E�M�UP��P�EjP�s����]��������������̸   �����������U��V�u��t���u6�EjP�s������u3�^]Ë��qt����t���t��U3�;P��I#�^]�����������P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������h~Ph^� �0������������������U��Vh~jh^� ���	�������t�@��t�M�UQRV�Ѓ�^]� 3�^]� �Vh~jh^� �����������t�@��tV�Ѓ�^�3�^���U��Vh~jh^� ����������t�@��t�M�UQRV�Ѓ�^]� ���^]� U���  Vh~jh^� ���S�������t/�@��t(�MWQ��x���VR�Ћ��E���b   ���_^��]� �u���c����N`�[������   �P�����   �E�����ݞ�  ��^��]� ����U��Vh~jh^� �����������t�@��t�M�UQRV�Ѓ�^]� ��������U��Vh~jh^� ����������t�@��t�M�UQ�MRQV�Ѓ�^]� ����U��Vh~j h^� ���I�������t�@ ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh~j$h^� �����������t�@$��t�MQV�Ѓ�^]� 3�^]� �����U��Vh~j(h^� ����������t�@(��t�M�UQ�MR�UQRV�Ѓ�^]� U��QVh~j,h^� ���x�������t �@,�E���t�E�MPQV�U���^��]� ��^��]� ��������U��Vh~j0h^� ���)�������t#�@0��t�E�M�U���$QRV�Ѓ�^]� 3�^]� ��������Vh~j4h^� �����������t�@4��tV�Ѓ�^�3�^���Vh~j8h^� ����������t�@8��tV�Ѓ�^�������U���`Vh~jDh^� ���v�������t(�@D��t!W�M�VQ�Ћ��E���   ���_^��]� �u��������^��]� ����U��Vh~jHh^� ����������t�@H��t
�MQV�Ѓ�^]� ������������U��Vh~jLh^� �����������t�@L��t�MQV�Ѓ�^]� ���^]� ����U��Vh~jPh^� ����������t�@P��t
�MQV�Ѓ�^]� ������������U��Vh~jTh^� ���Y�������t�@T��t
�MQV�Ѓ�^]� ������������U��Vh~jXh^� ����������t.�@X��t'�M �UQ�MR�UQ�MR�UQ�MRQV�Ѓ� ^]� 3�^]� �������������Vh~j`h^� ����������t�@`��tV�Ѓ�^�3�^���U��Vh~jdh^� ����������t�@d��t�MQV�Ѓ�^]� 3�^]� �����U���Vh~jhh^� ���F�������t1�@h��t*�MQ�U�VR�Ћu��P�������M�������^��]� �u�������^��]� �����������Vh~jph^� �����������t�@p��tV�Ѓ�^Ã��^��Vh~jlh^� ����������t�@l��tV�Ѓ�^Ã��^��Vh~jth^� ���|�������t�@t��tV�Ѓ�^�3�^���U��Vh~jxh^� ���I�������t�@x��t
�MQV�Ѓ�^]� ������������Vh~j|h^� ����������t�@|��tV�Ѓ�^�������Vh~h�   h^� �����������t���   ��tV�Ѓ�^�U��Vh~h�   h^� ����������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������U��Vh~h�   h^� ���V�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U���Vh~h�   h^� ����������tU���   ��tKW�M�VQ�Ћ�}�u���B�HV�ы�}�B�HVW�ы�}�B�P�M�Q�҃�_��^��]� ��}�H�u�QV�҃���^��]� ����������Vh~h�   h^� ���i�������t���   ��tV�Ѓ�^Ã��^������������U��Vh~h�   h^� ���&�������t���   ��t
�MQV�Ѓ�^]� ������U��Vh~h�   h^� �����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh~h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������Vh~h�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U��Vh~h�   h^� ����������t%���   ��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���U��Vh~h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ���^]� ����������U��Vh~h�   h^� ���f�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh~h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh~h�   h^� �����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh~h�   h^� ���v�������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������Vh~h�   h^� ���)�������t���   ��tV�Ѓ�^�3�^�������������Vh~h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������Vh~h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh~h�   h^� ���i�������t���   ��tV�Ѓ�^�3�^�������������U��Vh~h�   h^� ���&�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������Vh~h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U���Vh~h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh~h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh~h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U���Vh~h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh~h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh~h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U��Vh~h�   h^� ����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��QVh~h�   h^� ���E�������t#���   �E���t�E�MPQV�U���^��]� ��^��]� ��U��Vh~h�   h^� �����������t!���   ��t�E�M�U���$QRV�Ѓ�^]� ���������U��Vh~h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh~h�   h^� ���V�������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh~h   h^� ����������t��   ��t�MQV�Ѓ�^]� 3�^]� ���������������Vh~h  h^� ����������t��  ��tV�Ѓ�^�3�^�������������U���Vh~h  h^� ���s�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh~h  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh~h  h^� ���s�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U��Vh~h  h^� �����������t��  ��t
�MQV�Ѓ�^]� ������U��Vh~h  h^� ����������t��  ��t
�MQV�Ѓ�^]� ������U��Vh~h  h^� ���v�������t��  ��t
�MQV�Ѓ�^]� ������Vh~h   h^� ���9�������t��   ��tV�Ѓ�^�3�^�������������U��Vh~h$  h^� �����������t��$  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh~h(  h^� ����������t!��(  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh~h,  h^� ���V�������t��,  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh~h0  h^� ���	�������t��0  ��tV�Ѓ�^�3�^�������������U��Vh~h4  h^� �����������t��4  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh~h8  h^� ���v�������t��8  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh~h<  h^� ���&�������t��<  ��t�M�UQ�MRQV�Ѓ�^]� ��������������U��Vh~h@  h^� �����������t��@  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh~hD  h^� ����������t��D  ��tV�Ѓ�^�3�^�������������U��Vh~hH  h^� ���F�������t��H  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh~hL  h^� �����������t��L  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh~hP  h^� ����������t!��P  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��QVh~hT  h^� ���U�������t'��T  �E���t�E�M�UPQRV�U���^��]� ��^��]� ��������������U��Vh~hX  h^� �����������t%��X  ��t�E�M�U���$Q�MRQV�Ѓ�^]� �����U��Vh~j<h^� ����������t�@<��t�M�UQRV�Ѓ�^]� ��������U��Vh~j@h^� ���i�������t�@@��t�MQV�Ѓ�^]� 3�^]� �����h~Ph�� �0������������������h~jh�� ��������uË@����U��V�u�> t/h~jh�� ���������t��U�M�@R�Ѓ��    ^]���U��Vh~jh�� ����������t �@��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh~jh�� ���Y�������t�@��t�M�UQR����^]� ����������U��Vh~jh�� ����������t�@��t�M�UQR����^]� ����������U��Vh~jh�� �����������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh~j h�� ����������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh~j$h�� ���9�������t �@$��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh~j(h�� �����������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh~j,h�� ����������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  �����������U��Vh~j0h�� ���9�������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh~j4h�� �����������t5�@4��t.�M(�E �UQ�M���$R�UQ�MR�UQ�MRQ����^]�$ 3�^]�$ ������U��QVh~j8h�� ����������t�@8�E���t�E�MPQ���U�^��]� ��^��]� ����������U��Vh~j<h�� ���9�������t�@<��t�M�UQR����^]� ����������U��Vh~j@h�� �����������t�@@��t�M�UQR����^]� 3�^]� ���U��Vh~jHh�� ����������t�@H��t�M�UQR����^]� 3�^]� ���U��Vh~jDh�� ���y�������t�@D��t�M�UQR����^]� 3�^]� ���U��QVh~jLh�� ���8�������t#�@L�E���t�E�EP�����$�U�^��]� ��^��]� �����U��Vh~jPh�� �����������t�@P��t�M�UQR����^]� 3�^]� ���U��Vh~jTh�� ����������t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh~jXh�� ���Y�������t(�@X��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh~j\h�� ���	�������t(�@\��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��V��~ Wu h~jh�� ��������t�@�ЉF�~��t6h~jh�� ��������t�@��t�M�UVQ�MRQ����_^]� _3�^]� ��������������U��V��W�~��t+h~jh�� �1�������t�@��t�M�UQR���Ѓ~ t1h~jh�� � �������t�N�U�M�@R�Ѓ��F    _^]� ����������U��V��~ u h~jh�� ��������t�@�ЉF�v��t+h~jh�� ��������t�@��t�M�UQR����^]� �������������U��V�q��t@h~jh�� �D�������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ��������������U��V�q��t<h~j h�� ���������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��SV��~ Wu h~jh�� ��������t�@�ЉF�}�]�M�UWSQR���:  ��t�N��t�E�UWSPR����_^[]� _^3�[]� �U��V�q��t8h~j(h�� �$�������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� ������U��I��t)�E$�E�UP�E���\$�E�$R�UPR����]�  3�]�  �������U��V�q��t<h~j0h�� ��������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �������������U��V�u�F��F�����������������\{  ����������D�Ez��^�P�P�]��������������N�X�N^�X]���U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��u�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A �A�A(�A�������������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E����X�X]� ��̋�3ɉ�H�H�H�V��V����FP���3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  S�]���s  ��؋�U��M�U�>�U��@�����@�U��@�B�@�������@���@�   ;����U��p  �w�����  �w�������F�B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]؋�R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ʍU��R���[�[������E��KH��P�E�SL��H�щKP�P�ST�H�KX�P�����S\��z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����M��}������3�3����u��u�|+�A�����B�4�u�0u��u�p�����u�u�U�E;�}�Q���E����U��U��1���@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���@�D��KX�@�U�����]��C���@�K0���@�KH���C ��C�@�K8���@�KP���C(��C�C@�H���@3����KX���U��r  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������]��E�E����]���E����]��E׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���@�   �KXE)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� ����������h~Ph_� ��������������������h~jh_� ��������uË@����U��V�u�> t/h~jh_� ��������t��U�M�@R�Ѓ��    ^]���U��Vh~jh_� ���I�������t�@��t�MQ����^]� 3�^]� �������U��Vh~jh_� ���	�������t�@��t�MQ����^]� 3�^]� �������U��Vh~jh_� �����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh~jh_� ���y�������t�@��t�MQ����^]� 3�^]� �������U��Vh~j h_� ���9�������t�@ ��t�MQ����^]� 3�^]� �������U��Vh~j$h_� �����������t�@$��t�MQ����^]� 2�^]� �������Vh~j(h_� ����������t�@(��t��^��3�^������Vh~j,h_� ����������t�@,��t��^��3�^������U��Vh~j0h_� ���Y�������t�@0��t�MQ����^]� 3�^]� �������U��Vh~j4h_� ����������t�@4��t�M�UQR����^]� ���^]� ��Vh~j8h_� �����������t�@8��t��^��3�^������U��Vh~j<h_� ����������t�@<��t�MQ����^]� ��������������U��Vh~j@h_� ���i�������t�@@��t�MQ����^]� ��������������U��Vh~jDh_� ���)�������t�@D��t�MQ����^]� 3�^]� �������U��Vh~jHh_� �����������t�@H��t�MQ����^]� ��������������Vh~jLh_� ����������t�@L��t��^��3�^������Vh~jPh_� ���|�������t�@P��t��^��3�^������Vh~jTh_� ���L�������t�@T��t��^��^��������Vh~jXh_� ����������t�@X��t��^��^��������Vh~j\h_� �����������t�@\��t��^��^��������U��Vh~j`h_� ����������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh~jdh_� ���y�������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh~jhh_� ���9�������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh~jlh_� �����������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh~jph_� ����������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh~jth_� ���Y�������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh~jxh_� ����������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh~j|h_� �����������t�@|��t�MQ����^]� 3�^]� �������U��Vh~h�   h_� ����������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh~h�   h_� ���F�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh~h�   h_� �����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh~h�   h_� ����������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������m�������_�U�^��[�U����U��������������������d  ����������D�Ez���P�P���]� �������E�����E����X�M��X��]� �������U���@�`��A���E�    �����]����]��]��X��������]����]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P�����F�@��R�M��{����~���Q�M��i����v;�t�v��P�M��S����M����m��M�u�_^[�M�UQR�M�������]� ����������̋Q3���|�	��t��~�    t@����u��3���������U��QV�u;��}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��|+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~#V�1�d$ ���   @u	�����t@����u�^���̋QV3���~�	�d$ ����ШtF����u��^���������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%���;��E���}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$�H��E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��������3�����U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�����FP����3����F�F^��U��SV��WV�����^S�����E3����~�~;�t_��}�Q���   hh���jIP�у��;�t9�}��t;��}�B���   hh���    jNQ�҃����uV������_^3�[]� �E�~_�F^�   []� ����������U��SV��WV������^S������}3Ƀ��N�N;���   9��   �G;���   ��}�Q���  hh���jlP�у����t=� t@�G��t9��}�Jhh���    ���  jqR�Ѓ����u���-���_^3�[]� �O�N�G�Q��    R�F�QP�  �����t�N�WP��QPR�x  ��_^�   []� ���������U��SV��WV������~W�����3Ƀ��N�N9M��   �E;���   ��    ��}�H���  hh�h�   S�҃����t=�} tH�E��tA��}�Q���  hh���h�   P�у����u���2���_^3�[]� �U�V�,�F   ��}�H���  hh�h�   j�҃����t��E�M�F�PSPQ�q  �E����t!�V�?�W�RWP�U  ��_^�   []� ��M�_^�   []� ���U��Q�A�E� ��~LS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U�����u�_^[�E��Ћ�]� ���������U��S�]V��3�W�~���F�F�CV;C��   �$���W����3��F�F��}�Q���   hh�jIj�Ѓ������   ��}�Q���   hh�jNj�Ѓ����uV�������_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� ����W�z���3��F�F��}�B���   hh�jIj�у����t[��}�B���   hh�jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP��������^]� ����������U��U��t�M��t�E��tPRQ�PV  ��]�����������̡�}�H���   ��U���}�H���   V�u�R�Ѓ��    ^]����������̡�}�P���   Q�Ѓ�������������U���}�P�EPQ���   �у�]� ̡�}�H�������U���}�H�AV�u�R�Ѓ��    ^]��������������U���}�H�AV�u�R�Ѓ��    ^]��������������U���}�P��Vh�  Q���   �E�P�ы�}���   �Q8P�ҋ��}���   ��U�R�Ѓ���^��]��������������̡�}�P�BQ�Ѓ����������������U���}�P�EPQ�J\�у�]� ����U���}�P�EP�EP�EP�EP�EPQ���   �у�]� �U���}�P�EP�EP�EP�EPQ�JX�у�]� �������̡�}�P�B Q��Y�U���}�P�EP�EP�EP�EPQ���   �у�]� �����U���}�P�EP�EP�EPQ�J�у�]� ������������U���}�H��   ]��������������U���}�P�R$]�����������������U���}�P�EP�EP�EP�EPQ�J(�у�]� ��������U���}�P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U���}�P�EP�EP�EP�EPQ�J,�у�]� ��������U���}V��H�QWV�ҋ���}�H�QV�ҋ�}�Q�M�R4Q�MQ�MQOWHPj j V�҃�(_^]� ���������������U���}�P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U���}�P�EP�EPQ�J@�у�]� U���}�P�EPQ�JD�у�]� ���̡�}�P�BLQ�Ѓ���������������̡�}�P�BLQ�Ѓ���������������̡�}�P�BPQ�Ѓ����������������U���}�P�EPQ�JT�у�]� ����U���}�P�EPQ�JT�у�]� ����U���}�P�EP�EPQ���   �у�]� �������������U���}�P�E���   ��VP�EPQ�M�Q�ҋu�    �F    ��}���   j P�BV�Ћ�}���   �
�E�P�у� ��^��]� ������̡�}�P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡�}�H�������U���}�H�AV�u�R�Ѓ��    ^]��������������U���}�P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U���}�P�EPQ�J�у�]� ���̡�}�P�BQ��Y�U���}�P�EP�EPQ�J�у�]� U��VW���Ԝ���M�U�x@�EPQR��辜���H ���_^]� �U��VW��褜���M�U�xD�EPQR��莜���H ���_^]� �V���x����xH u3�^�W���f����΍xH�\����H �_^�����U��V���E����xL u3�^]� W���0����M�U�xL�EPQR�������H ���_^]� �������������U��V��������xP u���^]� W���ߛ���M�U�xP�EP�EQRP���ś���H ���_^]� ��������U��V��襛���xT u���^]� W��菛���M�xT�EPQ���}����H ���_^]� U���S�]VW���t.�M��vj�����O����xL�E�P���A����H ��ҍM��j���}��tZ��}�H�A�U�R�Ћ�}�Q�J�E�WP�ы�}�B�P�M�Q�҃��������@@��t��}�QWP�B�Ѓ�_^[��]� ������U��VW��贚���xH�EP��覚���H ���_^]� ���������U��VW��脚���M�U�xD�EP�EQRP���j����H ���_^]� �������������U��V���E����xP u
�����^]� W���-����M�U�xP�EP�EQ�MR�UPQR�������H ���_^]� ��������������U��V�������xT u
�����^]� W���͙���M�xT�EPQ��軙���H ���_^]� ��������������U��V��蕙���xX tW��臙���xX�EP���y����H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��  ����t.�E�;�t'��}�J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡�}�H��   ��U���}�H��$  V�u�R�Ѓ��    ^]�����������U���}�UV��H��(  VR�Ѓ���^]� �����������U���}�P�EQ��,  P�у�]� �U���}�P�EQ��,  P�у����@]� �����������̡�}�H��0  ���}�H��4  ��U��E��t�@�3���}�RP��8  Q�Ѓ�]� �����U���}�P�EPQ��<  �у�]� �U���}�P�EP�EP�EPQ��@  �у�]� ���������U���}�P�EP�EPQ��D  �у�]� �������������U���}�P�EPQ��H  �у�]� �U���}�P�E��L  ��VWPQ�M�Q�ҋu����}�H�QV�ҡ�}�H�QVW�ҡ�}�H�A�U�R�Ѓ�_��^��]� ��������������̡�}�P��T  Q�Ѓ������������̡�}�P��P  Q�Ѓ�������������U���}�P�EPQ��X  �у�]� ̡�}�H��\  ��U���}�H��`  V�u�R�Ѓ��    ^]�����������U���}�P�EP�EP�EP�EP�EPQ��d  �у�]� �U���}�P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w���2�����3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7���O����xP t$S���A���j j �XPj�FP���-����H ���[�    �~` t��}�H�V`�AR�Ѓ��F`    _^������������U��SV��Fx��}�Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR��������u#���h����}�H��0  h�   �҃��E�~P��������j j jW�N����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ��}�Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ������F|��u�E�~x��t�    �F`_^]� �M�Fx������t�3�_^]� U��QVW�}����	  ��}�H�QhV�҃�����}u"�H��0  h��h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���o  �EF;u�|�UR������_�   ^��]� �������������U��QVW�}�����  ��}�H�QhV�҃�����}u"�H��0  h��h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'����}�QP�Bh�Ѓ���t�M��R���  F;u�|ʍEP������_�   ^��]� �������������h��h�   h ~h�   �w�������t�������3��������V���(����N^��������������������U��VW�}�7��t��������N����V�]������    _^]�U���}�PH�EPQ���  �у�]� �U���}�P�B4VW�}j��h�  ���ЋMWQ���  _^]� ��������������U��V���PXW�ҋ}P����,�����Et�_�   ^]� �M�UPWQR���q  _^]� �����������U��S�]VW��j ���*���8�  �}uI�~ uC��}�P���   j h�  ���Ѕ�u��}�QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ���  _^[]� ��������U��EP�A    ��
����]� �����̸   �A� ������A   � ������U���@S�]VW����`��u�G   �}  ����   �M3�V�)���8�  u4����P�w�
����}�P�M�B4��jh�  ��_^�C�[��]� �MV�u)���8�  u�E�M��RPQ����_^�   [��]� �MV�E)���8�  t�MV�4)���8��  ��}�P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P�-���3��؃��u�;�t��}�QH���  VS�Ѓ��E��M�;O�f  9w�]  ��}�B�M���   Vh�  �҅�u!��}�P�M���   Vh�  �Ѕ��  ��}�Q�M�B4Vh�  ��;�t
V���������E��G��}���   ���   �Ћ]�E�;���   ;���   S�'���M���jQ�ˉu��uĉuȉủuЉu؉u�������U�E��ˉu��u�u�U�E��]��E�   �������t!��t��t�u���E�   ��E�   ��E�   �����M�;�t�>����BX�M�Q����P�����M܃�;�t�<���M��$���M��$���M��s���]�M�U�EQSRP���=  _^[��]� �M��\s��_^�   [��]� ��������������h~Ph�f �О�����������������U��h~jh�f 謞������t
�@��t]�����]�������U��Vh~jh�f �{���������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�j����E�NP�у�4�M��������^]ÍM�������^]��U��h~jh�f ��������t
�@��t]��3�]��������U��h~jh�f �ܝ������t�x t�P]��3�]������V��FW��u�~��N�<��u�< ��u_3�^á�}�H�F��  h�j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� }(�V;Vu��������t�F�N��    �F9~|؋V;Vu���������t��F�N�U���F_�   ^]� ��������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T����H;ǉ�F�M���F_�   ^]� ����U��E��|2�Q;�}+J;Q}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�s���3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�T��}���3����_�F�F^��������������U���SV�uW���^S�}��F���3���F�F�O�N�W���V9G�E~|��I �O���F�U�9FuL��u�~��~��t���< ��tY��}�H���  h�j8��    RP�у���t0�~�}���V��M����E�F@;G�E|�_^�   [��]� _^3�[��]� U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|���P�����_^]� �U����E�Qj�E��ARP�M��E�\�苿����]� �����U����Q�Ej�E��A�MRPQ�M��E�\�觿����]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q����t!�A��t�B�A�Q�P�A    �A    �̋�� d��@��HV3��q�q�P�r�r���p�p�p�P�H^������V���d������F3��F�;�t�N;�t�H�F�N�H�V�V�F�F�;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3���;�t�F;�t�A�F�N�H�V�V�Et	V�6�������^]� ������������U��V��W�~W�T������3����E��F�Ft	V�������_��^]� ������U��V��������Et	V���������^]� ��������������̸   � ��������� ������������̃��� ����������� �������������U���}�H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� ��}�Q0�F�M���   PQW�ҋF��^_]� U���}�H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U���}�H���  ]��������������U���}�H���  ]��������������U���}�P�EP�EP�EP�EPQ���   �у�]� �����U���}�E�P�EP�E���\$�E�$PQ���   �у�]� �������������U���}�P�EP�EP�EPQ���   �у�]� ��������̡�}�P���   Q�Ѓ�������������U���}�P�EP�EP�EPQ���   �у�]� ���������U���}�P�EP�EPQ���   �у�]� �������������U���}�H�U�ApR�Ѓ�]� �����U���}�P�EP�EPQ���  �у�]� �������������U���}�P�EP�EPQ���  �у�]� �������������U���}�P�EP�EPQ���  �у�]� �������������U���}�P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P�  ��R���E�P���ҡ�}�P�B<�M��Ћ}��t0j �M�QW�Qn������u��}�B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4���Т�E���E� '�E�`'�E��'�E��&�E�'�E��ǅx�����ǅ|���p��E�0'�E�p'�E��&�E�@'�E��'�E��&�E� '�E�P'�E� ��E����EĐ'�������}���B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۉ]���u��}�H�A�UR�Ѓ�^3�[��]Ë�}�Q�B<W�M3��Ѕ��'  �����E���tq�MQ�M��y���Wh���M������P�M��b����u�Wj��U�R�E�P��\���Q�_?������P��x���R������P�E�P������P��������E���t�E� �� t�M����耳����t��x�������m�����t��\�������Z�����t�M̃���J�����t��}�Q�J�E�P����у���t�M�� ����}� t"�U(�E$�M�R�UP�EQ�MRPQ���������U�R��������E$�M�UVP�Ej QRP�����������}�Q�J�EP�у���_^[��]����������������U��E�M�UP�EQ�Mj RPQ������]�������������̋�`<����������̋�`L����������̋�`0����������̋�`P����������̋�`����������̋�`$����������̋�`4����������̋�`D����������̋�`T����������̋�`(����������̋�`8����������̋�`H����������̋�`����������̋�`,��U���V�u��u��=  �@�E��=  ���E�F�}� �E�u�E�H�����   �� ��   S�]W�   ;�s��uS�7  Y��u�   �F�Xt}��u�]��}���6  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPW�u�j �O6  ��$��u������E�t	�M����_[^�Ë�U��V��<  �@�u��<  jh   �F�)=  YY�F��th   �86  P�v�,  ���F   ��6  �f �F��^]Ë�WhDf������uV�(~V��  �����~Y|�^��_�hDf����}V�(~V�  �����~Y|�^Ë�U��E��V��}k�(~P�  Y��^]� ���}k�(~P�  YË�U���u�d0  Y��t]�=  ]ËI�m����t�j���Ë�U��V��������EtV�����Y��^]� ��U��E���t�Bm����t�j���]Ë�U��Qj �M��@���h�~������%�~ Y�M��N����á�~Ë�U��=�~ uh*��~��  Y�E��~]�j�'��/>  j �M�������}�e� �w��GN���8 t��l����t�j�����w��w�>  �M��Y�M�������E>  Ë�U��Qj �M�������ȋ j��~�������~��u�M������Ë�U��=�~ uh�*����Yj�����Y��t��~��M�H�3���~]Ë�U��E�xP v�xTr�@@���@Pj � L  YY]�j�J��4=  ��u��F   3��E��F�F�F�Ehp��N�l��F��������c=  � j�x���<  ��u��l�V�E�   ����Yj j�N�����t��$=  Ë�U��V�������EtV�����Y��^]� j����<  ��~����u{P�M��2�����~!u�����uXj4����Y�ȉM��E���t
V�������3�V�E� ������N�F?   �$t�������Ή5�~�j����~��~�M���M���������i<  Ë�U��E�xVWr�p��pj j �J  YY��u����}P�O<�t�����tVj �wJ  YY��u�p�P�OX�T���_^]Ë�U��VW���w ��vW�u�V�6����u�_^]� ��U��V�uWj ��������F��t�8P����Y�ǅ�u�F �f ��t�8P�}���Y�ǅ�u�f  _^]Ë�U��V�u�~ v�F���~�F���~ V����Y�N$��tj�E���^]Ë�Vj���&���P��2  YY��^Ë�V���6�0  �6����YY^��1�.  Y��1�5  YË�U���V�u��u�7  �@�E��P7  ���E�F�}� �E�u�E�H�����   �� ��   S�]��   s!��uS�1  Y��u�   �F�X��   ��u�]��}��0  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPh   �u�j ��/  ��$��u������E�t	�M����[^�Ë�U��V�u���}��������^]� ����5�����U��V������"����EtV����Y��^]� jD����E9  h���M��%����e� �E�P�M�����hl?�E�P�  �jD����9  h���M�������e� �E�P�M��P���h<J�E�P��  ̋�U��V�u���>��������^]� ��U��USVW�ڋ�����   ��@t����t��3Ɂ�;���3�A;�t����@��u��������� u3��^��t%��t �uh���u�H  ����t	P�  Y���u���fV�u�`H  ������t���tjj V�.  ����tV�ŋ�_^[]Ë�U���  �Pg3ŉE��Eh  Ph  ������Pj �~K  ����t3���u�������uP��������M�3���  �Ë�U���u� �]Ë�U���u�$�]Ë�U���u�(�]Ë�U���u�,�]Ë�U���f��u]�#6  �MH��f��]����@��f��t����f��
r��̋L$WSV��|$��to�q��tU���L$���:�t��t���:�t
��u�^[_3�Ê��:�u�~��a��t(���:�u��A��t�f���:�t��3�^[_���J  �G�^[_Ë�^[_Ë�U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$����U��QQSVWd�5    �u��E�z2j �u�u��u�Z} �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�XV  �� �E�_^[�E���]Ë�U��V��u�N3��  j V�v�vj �u�v�u�V  �� ^]Ë�U���8S�}#  u��3�M�3�@�   �e� �E��3�Pg�M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E��2Y  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M�  �E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u��T  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����-���u�[  �M�N��k���M9H};H~���u	�M�]�u�} }ʋEF�0�E�;_w;�v�t[  ��k�E�_^[�Ë�U��EV�u���W  ���   �F�W  ���   ��^]Ë�U���W  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V�yW  �u;��   u�iW  �N���   ^]��XW  ���   �	�H;�t���x u�^]��Z  �N�H�ҋ�U����Pg�e� �M�3��M�E��E�E�E@�E��2�M��E�d�    �E�E�d�    �uQ�u��Z  �ȋE�d�    ����;Pgu����Z  ��Q�D���[  YË�U��V��������EtV����Y��^]� ��U��E��	Q��	P�/\  ��Y�Y@]� ��U��E��t���8��  uP�  Y]Ë�U��EV���F ��uc�:V  �F�Hl��Hh�N�;Xnt�pm�Hpu�I5  ��F;xlt�F�pm�Hpu�R^  �F�F�@pu�Hp�F�
���@�F��^]� ��U����Pg3ŉE�S3�V;�u�(c  j^SSSSS�0�P  ���5  �uW�b  YY;Er��ЋU��H;�u ��8t�<a|<z, �A8u�3���   j�p�   SSj�WVQR�O'  �ȃ�$�M�;�u�b  � *   �b  � �   9Ms��b  j"�^���;�~Ej�3�X���r9�A=   w�b  ��;�t� ��  �P��  Y;�t	� ��  ���M�E���]�9]�u�.b  �    냋U�j�pQ�u�j�WV�pR�&  ��$��t�u��uW��   �������a  j*Y����u������Y�ƍe�^[�M�3��}����Ë�U���W�u�M�������}�E�P�u�_����}� YY_t�M��ap��Ë�U��j �u�u������]Ë�U��S3�9luA�E;�u�aa  SSSSS�    �	  ��3��/��8t)�
��a|
��z�� �
B8u��Sj��u�X����E��[]Ë�U��MS3�VW;�t�};�w��`  j^�0SSSSS�#	  �����0�u;�u��ڋъ�BF:�tOu�;�u���`  j"Y�����3�_^[]������̋T$�L$��ti3��D$��u��   r�=�� t�Wa  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$ø)���o��o���oĝ��o����of���o��o����o��� p��pq�Ë�U�������Mm  �} �Ht��l  ��]����U��WV�u�M�}�����;�v;���  ��   r�=�� tWV����;�^_u^_]�m  ��   u������r*��$�<��Ǻ   ��r����$�(;�$�$<��$��;�8;d;�;#ъ��F�G�F���G������r���$�<�I #ъ��F���G������r���$�<�#ъ���������r���$�<�I <�;�;�;�;�;�;�;�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�<��$<,<8<L<�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��=�����$�`=�I �Ǻ   ��r��+��$��<�$��=��<�<=�F#шG��������r�����$��=�I �F#шG�F���G������r�����$��=��F#шG�F�G�F���G�������V�������$��=�I d=l=t=|=�=�=�=�=�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��=���=�=�=�=�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ���` �` � X�Ë�U��S�]VW���X����t&P�|(  ��FV�=  YY�G��t�3VP��������g �G   ��_^[]� ��U��S�]V���X��C�F���CWt1��t'P�(  ��GW��  YY�F��t�sWP�D������	�f ��F_��^[]� �y �X�t	�q��  YËA��u�`�Ë�U��V�EP�������x���^]� ��U��V�u���R����x���^]� �x�������U��V�������EtV�i���Y��^]� ��U��V���x��c����EtV�B���Y��^]� ��U��V�uW3�;�u3��e9}u�vZ  j^�0WWWWW�  �����E9}t9urV�u�u�  �����uW�u������9}t�9us�'Z  j"Y����jX_^]�������������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[Ë�U��EVW3�;�tG9}u�CY  j^�0WWWWW�k  �����)9}t�9Es�Y  j"Y�����P�u�u�_�����3�_^]Ë�U��E�L]Ë�U���(  �Pg3ŉE������� SjL������j P������������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������D�j ���@���(���P�<���u��uj�g  Yh ��8�P�4��M�3�[�}����Ë�U���5L��G  Y��t]��j��f  Y]����3�PPPPP�������Ë�U��� �EVWjY����}��E��E_�E�^��t� t�E� @��E�P�u��u��u��H��� jhxJ�ys  �u��tu�=|�uCj�kh  Y�e� V�h  Y�E��t	VP�h  YY�E������   �}� u7�u�
j�Wg  Y�Vj �5���P���u��V  ���L�P�V  �Y�=s  �jh�J��r  3��}�3��u;���;�u �V  �    WWWWW����������   V�}u  Y�}��F@uwV�z  Y���t���t�����ȃ����@����s�A$u)���t���t���������@����s�@$�t�
V  �    WWWWW�1������M��9}�u�Nx
��A��V��u  Y�E��E������   �E��Dr  ËuV�3u  Y�jh�J��q  3��}�3��u;���;�u �U  �    WWWWW����������   V�yt  Y�}��F@uwV�y  Y���t���t�����ȃ����@����s�A$u)���t���t���������@����s�@$�t�U  �    WWWWW�-������M��9}�u!�Nx��E�����V�u�x  YY�E��E������   �E��8q  ËuV�'t  YË�U��V�u�F@WuyV�Gx  Y��s���t���t�ȃ��������@�����A$u&���t���t�ȃ������@�����@$�t�:T  3�WWWWW�    �_���������JS�]���t=�F�u��y2�u.3�9~uV�Ey  Y�;Fu9~u@���F@�t8t@����[_^]È�F�F�����F��%�   ��jh�J��o  3�3�9u��;�u�S  �    VVVVV�����������+�u�r  Y�u��u�u�����YY�E��E������	   �E���o  ��u��r  YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV��v  YP��  ��;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�]v  P�E�  Y��Y��3�^]�jh�J��n  3��}�}�j��c  Y�}�3��u�;5`���   �@���98t^� �@�tVPV�q  YY3�B�U��@����H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u�@��4�V�q  YY��E������   �}�E�t�E��In  �j�+b  Y�jh K��m  3�9uu	V����Y�'�u�p  Y�u��u����Y�E��E������	   �E���m  ��u��p  Y�j�����Y�jh@K�m  3ۉ]�3��u;���;�u �<Q  �    SSSSS�c���������   �E��t	;�t��@u�;�t��@u�}�G�=���v뷋}����uV��o  Y�]�V����V�\  YY�f�����N�Et���Fj_�-�E;�u W�"  Y;�u�L��M����N  �	��   �N�~�F��^�E������	   �E���l  ��u��o  YË�U���SVW3�9}t$9}t�u;�u�?P  WWWWW�    �f�����3�_^[�ËM;�tڃ��3��u9Ew͋}�}�F  �M��}��t�F�E���E�   ����   �N��  t/�F��t(��   ��;�r��W�u��6��
  )~>��+�}��O;]�rO��tV�S���Y��u}�}� ��t	3ҋ��u�+�W�u�V�-s  YP�8|  �����ta��;�w��M�+�;�rP�}��)�E�� VP�-s  YY���t)�E��FK�E����E�   ���A����E������N ��+�3��u������N �E���jh`K�2k  3�9ut)9ut$3�9u��;�u ��N  �    VVVVV�������3��@k  ��u�m  Y�u��u�u�u�u�=������E��E������   �E����u��m  YË�U��W3�9}u�lN  WWWWW�    ����������AV�u;�u�GN  WWWWW�    �n����������u�'�  Y�ȉ#ʃ���V;�t3�^_]Ë�U��V�u�F��u��M  �    ����g���}�FuV�y�  E�e YV�����FY��y����F��t�t�   u�F   �u�uV�Rq  YP�V�  3Ƀ������I��^]�jh�K�i  3�3�9u��;�u�gM  �    VVVVV����������>�};�t
��t��u��u�?l  Y�u�W�u�u�������E��E������	   �E��i  ��u�l  YË�U��V3�9uu��L  VVVVV�    �����������E;�t�V�p�0�u薂  ��^]Ë�U��SV�uW3����;�u�L  WWWWW�    ���������B�F�t7V�:���V����z  V�&p  P�+�  ����}�����F;�t
P����Y�~�~��_^[]�jh�K�wh  �M��3��u3�;���;�u� L  �    WWWWW�G����������F@t�~�E��zh  �V��j  Y�}�V�*���Y�E��E������   �ՋuV�Gk  YË�U���u�T���u�L��3���tP��K  Y���]�3�]Ë�U��� WV�0  3�Y;�u�~K  WWWWW�    ����������49}t޹����E�I   �u�u��M�;�w�E��u�E��u�uP�U��_�Ë�U��V�u�EPj �uh���z�����^]Ë�U��Q�e� S�]��u3��   W��ru�{���vn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9}�r��?�@��I��F�@��I��<�@��I��2�@��I��(�M�E����t:u@A�E�9]�r�3�_[��� �	+����U��j
j �u�~�  ��]��5l��d:  Y��t��j苔  jj �]  ���>  ��U��EVW��u|P�Y  Y��u3��  �">  ��u�5Y  ���3�  �\������  �T��j  ��}�:  ����  ��| 薚  ��|j �g�  Y��u�P�   ��l  ��3�;�u19=P~��P9=��u���  9}u{�l  �9:  �X  �j��uY��9  h  j��  ��YY;��6���V�54h�5x�O9  Y�Ѕ�tWV�-:  YY�X��N���V����Y�������uW�<  Y3�@_^]� jh�K�
e  ����]3�@�E��u9P��   �e� ;�t��u.�����tWVS�ЉE�}� ��   WVS�r����E����   WVS�ra���E��u$��u WPS�^a��Wj S�B��������tWj S�Ѕ�t��u&WVS�"�����u!E�}� t�����tWVS�ЉE��E������E���E��	PQ� �  YYËe��E�����3��fd  Ë�U��}u���  �u�M�U�����Y]� ����̃=� �0�  ���\$�D$%�  =�  u�<$f�$f��f���d$���  � �~D$f(��f(�f(�fs�4f~�fT��f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$连  ���D$��~D$f��f(�f��=�  |!=2  �fT���\�f�L$�D$����f���fV��fT��f�\$�D$���������������̃=�� t-U�������$�,$�Ã=�� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$��jh�K�b  �e� �u;5l�w"j�W  Y�e� V�_  Y�E��E������	   �E��b  �j��U  YË�U��V�u�����   SW�=`��=�� u耑  j�Ώ  h�   躓  YY�|���u��t���3�@P���uV�S���Y��u��uF�����Vj �5���׋؅�u.j^9��t�u�e�  Y��t�u�{�����D  �0��D  �0_��[�V�>�  Y��D  �    3�^]�������������U��WV�u�M�}�����;�v;���  ��   r�=�� tWV����;�^_u^_]�R  ��   u������r*��$�W��Ǻ   ��r����$�V�$�W��$��V�(VTVxV#ъ��F�G�F���G������r���$�W�I #ъ��F���G������r���$�W�#ъ���������r���$�W�I �V�V�V�V�V�V�V�V�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�W��WW(W<W�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��X�����$�PX�I �Ǻ   ��r��+��$��W�$��X��W�W X�F#шG��������r�����$��X�I �F#шG�F���G������r�����$��X��F#шG�F�G�F���G�������V�������$��X�I TX\XdXlXtX|X�X�X�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��X���X�X�X�X�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U��QSVW�5��y1  �5����}��i1  ��YY;���   ��+ߍC��rwW�r�  ���CY;�sH�   ;�s���;�rP�u���  YY��u�G;�r@P�u���  YY��t1��P�4��0  Y���u�v0  ���V�k0  Y���EY�3�_^[�Ë�Vjj �G  ��V�D0  ��������ujX^Ã& 3�^�jh L�\  �Ԏ  �e� �u�����Y�E��E������	   �E��\  �賎  Ë�U���u���������YH]�������������̺�g遝  ��g���  �Ƀ=Ht����D�  �����z�����������������̃��$药  �   ��ÍT$�8�  R��<$�D$tQf�<$t��  �   �u���=D �c�  �   ��g�`�  �  �u,��� u%�|$ u���Ů  �"��� u�|$ u�%   �t����-�t�   �=D ��  �   ��g��  ZË�U����Pg3ŉE�SV3�W��9du8SS3�GWh �h   S�p���t�=d��L���xu
�d   9]~"�M�EI8t@;�u�����E+�H;E}@�E�d����  ;���  ����  �]�9] u��@�E �5l�3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�l>  ��;�t� ��  �P�r���Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5p�SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�=  ��;�tj���  ���P����Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�p���t"SS9]uSS��u�u�u�VS�u �h��E�V�����Y�u�������E�Y�Y  �]�]�9]u��@�E9] u��@�E �u耭  Y�E���u3��!  ;E ��   SS�MQ�uP�u 螭  ���E�;�tԋ5d�SS�uP�u�u�։E�;�u3��   ~=���w8��=   w�<  ��;�t����  ���P����Y;�t	� ��  �����3�;�t��u�SW�^������u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u���  ���u������#u�W�����Y��u�u�u�u�u�u�d���9]�t	�u��L���Y�E�;�t9EtP�9���Y�ƍe�_^[�M�3������Ë�U����u�M������u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap����-  �ȋAl;Xnt�pm�Qpu�  ���   Ë�U����u�M������E����   ~�E�Pj�u蟭  ������   �M�H���}� t�M��ap��Ë�U��=l u�E�Hn�A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u� �  ������   �M�H���}� t�M��ap��Ë�U��=l u�E�Hn�A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u衬  ������   �M�H���}� t�M��ap��Ë�U��=l u�E�Hn�A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Ph�   �u��  ������   �M�H%�   �}� t�M��ap��Ë�U��=l u�E�Hn�A%�   ]�j �u�~���YY]Ë�U����u�M������E����   ~�E�Pj�u蜫  ������   �M�H���}� t�M��ap��Ë�U��=l u�E�Hn�A��]�j �u����YY]Ë�U���L�Pg3ŉE�S3�V�uW�]ԉ]�]��]؉]܉u��]�9^�  �F9u P�F0h  P�E�SP�x�  ������  j�  j��  W�E��  jW�E��  jW�E��  jh  �E��  ��$�E�9]��|  9]��s  ;��k  9]��b  9]��Y  �Eԉ3��M܈@=   |�E�P�v�t����/  �}��%  �E���E�~-8]�t(�E�:�t�x�����M�� �G;�~�@@8X�uۋE�SS�v   Ph   �u܉E�jS�a�  �� ����  �M��E�S�v��   W���   QW@Ph   �vS������$����  �E�S�v�   WP�E�W@Ph   �vS�U�����$���`  �E�}����   3҃}�f��U؉Mč��   �_�Z��M����   �MȈ~S8]�tN�M�M�:�tB�I���;ʉM�'��H   ��M��E� �  f�AA�M̋M��	9M�~�M�AA�M�8Y�u�h�   ��   QP�]���j��   PW�N����E�j��   QP�<������   ��$;�tKP����u@���   -�   P�������   ��   +�P�s������   +�P�e������   �Z������E��    ���   �E����   �Eĉ��   �E����   �Eȉ��   �EЉ��   �u�����Y���m�u������u�������u�������u������3ۃ�C�ˍ��   �;�tP������   ǆ�   �ǆ�   ��ǆ�   �ǆ�      3��M�_^3�[�������X'  �ȋAl;Xnt�pm�Qpu�r  �@��2'  �ȋAl;Xnt�pm�Qpu�L  ��Ë�U��VW3��u�������Y��u'9hvV�����  ;hv��������uʋ�_^]Ë�U��VW3�j �u�u赩  ������u'9hvV�����  ;hv��������uË�_^]Ë�U��VW3��u�u艪  ��YY��u,9Et'9hvV�����  ;hv��������u���_^]Ë�U��VW3��u�u�u�S�  ������u,9Et'9hvV�����  ;hv��������u���_^]��̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U���(  �Pg3ŉE�� hVtj
�}  Y�/�  ��tj�1�  Y� h��   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P�V�������������(�����0���j ǅ����  @��������,����@���(���P�<�j�8�  ̋�U��M� h�U#U��#�ʉ h]�Pd�5    �D$+d$SVW�(��Pg3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(��Pg3�P�e��u��E������E�d�    ËM�d�    Y__^[��]QË�U��SV�u���   3�W;�to=wth���   ;�t^9uZ���   ;�t9uP�������   �P�  YY���   ;�t9uP�r������   � �  YY���   �Z������   �O���YY���   ;�tD9u@���   -�   P�.������   ��   +�P�������   +�P�������   ���������   �=Pvt9��   uP药  �7�����YY�~P�E   ��xmt�;�t9uP����Y9_�t�G;�t9uP����Y���Mu�V����Y_^[]Ë�U��SV�5�W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�xmt	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5�W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�xmt	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�V���t��t;�tWj6Y���  P����Y_^Å�t7��t3V�0;�t(W�8����Y��tV�����> Yu���mtV�3���Y��^�3��jh L�wJ  �   ��pm�Fpt"�~l t�   �pl��uj �|  Y���J  �j�F?  Y�e� �Fl�=Xn�i����E��E������   ��j�A>  Y�u�áXn�H���H�����   �\n���   �w���   �@w���   ��g���   �DwË�U��SW�}3�;�~,V�u���6�u�u�0�  ����tSSSSS�V�����Ou�^_[]Ë�U��SVW�}h�   3�SW�y����u�����u3���   <.u4�F8t-jP���   jP萴  ����tSSSSS����������   ��h�V�]� �  ;��   �} �<0�u��@��   ��.��   PVj@�u�;�}u��@sw��_trP�EVj@��@��}u`��s[��t��,uRP�EVj��P���  ����t3�PPPPP�Y�������,�'����������E�wh�V�{�  ��YY�X������_^[]Ë�U��SV�uV�u�u�������3ۅ�tSSSSS��������F@8tPh�j�u�u�Q��������   8^[tPh��j�u�u�/�����]Ë�U���S3�ChU  �]�� ���Y�E���U  W�x� ��]��^�CH�0�E�h$��5\�jhQ  W������E���E��E�\�h �hQ  W�
�  ����t3�PPPPP�.������sX�E��0�E#  YY��t�e� �E��E��E����0�CH�0�E�E�h$��0jhQ  W�Z������}���|��}� uI�FP����tP�Ӆ�u	�vP�a���Y�FT��tP�Ӆ�u	�vT�J���Y�E�fT �fL �FP�~H���N�u��,����FP�=�3�Y;�tP�ׅ�u	�vP����Y�FT;�tP�ׅ�u	�vT�����Y�Fh�^T�^L�^P�^H_[�Ë�U���   �Pg3ŉE��ESV�uW�}��d����E��\�����`����r  �   �H(��T����H,�X �   ��X�����h�������  ��d��� ��  �} ��  �>CuW�~ uQht��u��d����t�����3���tVVVVV������;�t3�f�f�Gf�G��`���;�t�0��d����G  V�������   Y��P���;�s,V��h����b!  YY����   V��X����L!  YY����   ��L��� ��l���VP����YY����   ��l���PSP��  ������   �C��T������l���PW��h����������> t
��P���;�r��L������@PVW��X����&�  ����t3�VVVVV�������3�9�\���tjS��\���������9�`���tj��T�����`�����������h����u��d�����������tVVVVV�#�������h����3��M�_^3�[�����Ë�U����  �Pg3ŉE�SW���^  �u����h���P��P���Ph�   ��x���PS���  ��������u3��  �E���0�sH��x���P�  YY���x  ��x���P������P��t��������YY��p�����t��CH�M��\����D���k���l���� ��X����1jP��d�����<���P�b����F��x���Q��t�����L�����p��������QP���������t3�PPPPP���������p�����l������CH��P����j��P���P��d�����������}��   ��h�����t��� �F�G$�O ��d����ǋV;t6���t������d�����D����P�H��D�������t�����d���|��"��t�����t�ǋ��P�W���d����H��t���uhj�v��x����vPjh��jj �=�  �� ��t93���  f!�Ex���@��r�h�   �5h��x���P�Ƶ  �����@�G��g �F��G���   �}u	��h����F�Ek�V��X�Y��t1��\�����p����CH�.�����X���Y��l������L����F������\���xmt-�E�����<0�7����u�7������sT������cL YY�M��p��������    �1�CH�M�_3�[�����Ë�U���   �Pg3ŉE��ESV3ۋ�W��h���;�t;�tP�����Y��  ���D0H��  ǅp���   ��t���;���  �9L�0  �yC�&  �y_�  ��h(�W���  ��YY����   +ǉ�p�����   �;;��   ǅl���   �\����p���PW�6��������u�6�����Y9�p���t��l���������~�Ch �S�N�  ��3�YY;�u	�;;��   ��l���QWS��x���h�   P�e�  ����tVVVVV���������l�����h�����x���Ƅ=x��� ����Y��t��t�����? t
G�? � ���3�9�t�����   ��h����u3��vSSSh�   ��x���PQ�"�����;�tZ�~H��t3�7��x���P�e  YY��tS��x����%���Y��u!�p������t���C����~�3�9�p���u9�t���t�D����M�_^3�[菾����jh@L�?  3ۉ]��}v�"  �    SSSSS�������3��,  �$  ���u��Q����Np�]�jh�   �;���YY���}�;���   j�3  Y�E�   �Nl�������]��   �u�M���P���Y�E�;���   9]thxm�u�^  YY��t
�l   j�X3  Y�E�   �^l���|���W����Y�Fpu2�pmu)�;�Xn�Z���j�Xn��PhЂ������������e� �   �-�}܋u�3�j�2  YËu�j�2  Y��W�N���W�p���YY�E������   �E���=  Ëu�fp��jhxL�=  3��u�3��];���;�u�G!  �    VVVVV�n�����3��{3��};���;�t�3�f97��;�t���  �E;�u�!  �    �ɉu�f93u ��   �    j��E�PhPg��  ���P�uWS��  ���E��E������	   �E��3=  ��u�#@  YË�U���SV�u3ۉ]�;�t9]u3��{  v3�f�W�};�u�o   SSSSS�    �������<  �u�M��~����E�;���   9XuH9]v�M��9f�f�8tAFF�M�;Mr�8]�t�E�`p��E���   8]�t�E�`p�����   �uVj�W�=l�j	�p��;���   �L���zt��  � *   3�f��   �E�u�E�;�t'��M�:�t�M���QP��  YY��tF8t!F9]�u��u+u�u�E�V�uj�p��;�uT�d  �M� *   3�f��-9Xu	W�����Y�1SSj�Wj	�p�l�;�u�-  � *   8]�t�E�`p�����H8]�t�M�ap�_^[�Ë�U���SV�u3ۉ]�;�u9]t*�9]w��  j^SSSSS�0����������   3�f�W�};�t��u�M��ܺ���E;Ev�E=���v	�  j�P�M�QP�uV����������u;�t3�f��k  � 8]�tk�M�ap��b@;�tH;Ev<�}�t,3�f��A  j"^SSSSS�0�i�����8]�t�E�`p����&�E�E�P   3�f�LF�;�t�8]�t�E�`p��E�_^[�Ë�U��j �u�u�u�u�u�������]����������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[Ë�U��V�EP��������4���^]� �4�������U��V���4��{����EtV�Z|��Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR�  YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =MOC�t=csm�u+�  ���    ��  �  ���    ~�  �   �3�]�jh�L�68  �}�]��   �s��s�u��\  �   � �e� ;ute���~;w|��  �����Oȋ1�u��E�   �y t�sh  S�O�t��  �e� ��u��-���YËe�e� �}�]�u��u���E������   ;ut�a  �s��7  Ë]�u��  ���    ~�  �   �Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�q  3�A��  ���3��jh�L�7  �M��t*�9csm�u"�A��t�@��t�e� P�q覲���E������7  �3�8E��Ëe��R  ̋�U��M�V�uƃy |�Q�I�42���^]Ë�U�����u
�c  �  �e� �? �E� ~SSV�E�@�@��p��~3�E����E�M�q�P�GE�P�_�������u
K�������E��E��E�;|�^[�E���j����u����X  ���    t��  �e� �  �M���|  �3  �Mj j ���   �
����j,h8M��5  �ً}�u�]�e� �G��E��v�E�P����YY�E���  ���   �E���  ���   �E���  ���   ��  �M���   �e� 3�@�E�E��u�uS�uW�j������E�e� �o�E������Ëe��  ��   �u�}�~�   �O��O�^�e� �E�;Fsk�ËP;�~@;H;�F�L�QVj W�������e� �e� �u�E������E    �   �E��5  ��E�맋}�u�E܉G��u��h���Y��
  �Mԉ��   ��
  �MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v����Y��t�uV�%���YY�jh`M�24  3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w���  YY����   SV���  YY����   �G��M��QP�����YY���   �}�E�p�tH��  YY����   SV��  YY����   �w�E�pV膷�������   ���t|��W�9Wu8�]�  YY��taSV�P�  YY��tT�w��W�E�p�_���YYPV�5������9�%�  YY��t)SV��  YY��t�w�
�  Y��t�j X��@�E���  �E������E��3�@Ëe��Q  3��3  �jh�M�2  �E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS�!�����FP�w����YYP�vS�����E������2  �3�@Ëe��  ̋�U��} t�uSV�u�V������}  �uuV��u �ŭ���7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP�O���]Ë�U��QQV�u�>  ���   W��  ���    t?��  ���   �z  9t+�>MOC�t#�u$�u �u�u�u�uV����������   �}� u�"  �u�E�P�E�PV�u W�1������E���;E�s[S;7|G;wB�G�O����H��t�y u*�X��@u"�u$�u�u j �u�u�u�u�����u���E��E���;E�r�[_^�Ë�U���,�MS�]�C=�   VW�E� �I��I����M�|;�|�h
  �u�csm�9>��  �~� ��  �F;�t=!�t="���   �~ ��   �  ���    ��  �  ���   �u�q  ���   jV�E�,�  YY��u��	  9>u&�~u �F;�t=!�t="�u�~ u�	  �&  ���    t|�  ���   �  �u3����   ����Y��uO3�9~�G�Lhh�O�����uF��;7|��	  j�u�d���YYh<��M��7���h�M�E�P蒻���u�csm�9>��  �~�~  �F;�t=!�t="��e  �}� ��   �E�P�E�P�u��u W�	��������E�;E���   �E�9��   ;G|�G�E�G�E��~l�F�@�X� �E��~#�v�P�u�E����������u�M��9E���M�E��}� ��(�u$�]��u �E��u��u�u�uV�u�K����u���E����]����}�} t
jV�:���YY�}� ��   �%���=!���   �����   V����Y����   �_  �Z  �U  ���   �J  �}$ �M���   Vu�u��u$让���uj�V�u�u�������v�����]�{ v&�} �)����u$�u �u�S�u�u�uV������� ��  ���    t�_  _^[�Ë�U��V�u��蔵���4���^]� ��U��SVW�  ��   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������� 3�@_^[]Ë�U��V�58h�5���օ�t!�4h���tP�58h���Ѕ�t���  �'�\�V�x���uV��]  Y��thL�P�|���t�u�ЉE�E^]�j ����YË�U��V�58h�5���օ�t!�4h���tP�58h���Ѕ�t���  �'�\�V�x���uV�X]  Y��thx�P�|���t�u�ЉE�E^]����� ��V�58h�������u�5t�e���Y��V�58h�����^á4h���tP�5|�;���Y�Ѓ4h��8h���tP����8h���  jh�M�+  �\�V�x���uV�\  Y�E�u�F\�3�G�~��t$hL�P�|��Ӊ��  hx��u��Ӊ��  �~pƆ�   CƆK  C�FhPhj�  Y�e� �vh���E������>   j�  Y�}��E�Fl��u�Xn�Fl�vl�O���Y�E������   �*  �3�G�uj�m  Y�j�d  YË�VW�L��54h�������Ћ���uNh  j������YY��t:V�54h�5x�����Y�Ѕ�tj V�����YY�X��N���	V�D���Y3�W���_��^Ë�V��������uj�v[  Y��^�jh N�)  �u����   �F$��tP�����Y�F,��tP����Y�F4��tP�۵��Y�F<��tP�͵��Y�F@��tP迵��Y�FD��tP豵��Y�FH��tP裵��Y�F\=�tP蒵��Yj�  Y�e� �~h��tW����u��PhtW�e���Y�E������W   j��  Y�E�   �~l��t#W�A���Y;=Xnt���mt�? uW�M���Y�E������   V����Y��(  � �uj�  YËuj�  YË�U��=4h�tK�} u'V�58h�5���օ�t�54h�58h���ЉE^j �54h�5x����Y���u�x����8h���t	j P���]Ë�VW�\�V�x���uV�Y  Y�����^  �5|�h��W��h��W�p��h��W�t��h��W�x�փ=p �5���|t�=t t�=x t��u$����t����p��5x�|����8h�����   �5tP�օ���   �[  �5p�����5t�p�����5x�t�����5|�x�u������|�v  ��teh��5p�����Y�У4h���tHh  j�6�����YY��t4V�54h�5x����Y�Ѕ�tj V�y���YY�X��N��3�@��$���3�_^�jh(N�j&  �����@x��t�e� ���3�@Ëe��E������6����&  ��~����@|��t������jhHN�&  �5�����Y��t�e� ���3�@Ëe��E������}����h��g���Y������������U���SQ�E���E��EU�u�M�m���  VW��_^��]�MU���   u�   Q�ö  ]Y[�� ��U���(  �������������5���=|�f���f���f�x�f�t�f�%p�f�-l������E ����E����E�����������  �������	 ���   �Pg�������Tg�������D���j�  Yj �@�h���<��=� uj�|  Yh	 ��8�P�4���jhhN�z$  j�|  Y�e� �u�N��t/�������E��t9u,�H�JP辰��Y�v走��Y�f �E������
   �i$  Ë���j�G  Y��������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�R���3��ȋ��~�~�~����~����Ph���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �Pg3ŉE�SW������P�v�t��   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R菥����C�C��u�j �v�������vPW������Pjj �O{  3�S�v������WPW������PW�vS������DS�v������WPW������Ph   �vS�^�����$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[�Р����jh�N�N!  �������pm�Gpt�l t�wh��uj ��R  Y���f!  �j�"  Y�e� �wh�u�;5xlt6��tV����u��PhtV�d���Y�xl�Gh�5xl�u�V���E������   뎋u�j��  YË�U���S3�S�M�薠��������u���   ���8]�tE�M��ap��<���u���   ����ۃ��u�E��@���   ��8]�t�E��`p���[�Ë�U��� �Pg3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9��l��   �E��0=�   r����  �p  ����  �d  ��P������R  �E�PW�t����3  h  �CVP询��3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�h����M��k�0�u����l�u��*�F��t(�>����E���|lD;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C���lZf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95���X�������M�_^3�[�˝����jh�N�I  �M���������}�������_h�u�u����E;C�W  h   �J���Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh����u�Fh=PhtP�@���Y�^hS�=����Fp��   �pm��   j�  Y�e� �C�Ă�C�Ȃ�C�̂3��E��}f�LCf�E��@��3��E�=  }�L��pj@��3��E�=   }��  ��xk@���5xl����u�xl=PhtP臩��Y�xlS���E������   �0j�  Y��%���u ��PhtS�Q���Y�   �    ��e� �E��  Ã= � uj��V���Y� �   3�Ë�U��3�9Ev�M�9 t@A;Er�]Ë�U��E3�;�hntA��-r�H��wjX]Ë�ln]�D���jY;��#���]�������u��oÃ���������u��oÃ�Ë�U��V������MQ�����Y�������0^]��������������Q�L$+ȃ����Y�:�  Q�L$+ȃ����Y�$�  U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh�N��  �e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E���  Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[���������3�Ë�U���V�u�M�������u�P�Ѭ  ��e�F�P�������Yu��P贬  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�脙���E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P��  �M��E��M��H��EP��  �E�M����Ë�U��j �u�u�u������]Ë�V����tV����@PV�V訜����^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M����A���3�;�u+����j_VVVVV�8�,������}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�����j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h��SV�)�����3ۅ�tSSSSS�=������N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F��t�90uj�APQ�%������}� t�E��`p�3�_^[�Ë�U���,�Pg3ŉE��ESVW�}j^V�M�Q�M�Q�p�0蒬  3ۃ�;�u�y���SSSSS�0褢�������o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q诪  ��;�t���u�E�SP�u��V�u��������M�_^3�[蜕���Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �Օ��9}}�}�u;�u+����j^WWWWW�0跡�����}� t�E�`p����  9}vЋE��� 9Ew	�Q���j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV蕦  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� �]�  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �	�  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V葖����u�E�8 u���} �4����$�p���WF蕪  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP�p�  0�F�U�����;�u��|��drj jdRP�J�  0��U�F����;�u��|��
rj j
RP�$�  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N�i�����u-�.���j^�03�PPPPP�T������}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V�˔�����}� t�E��`p�3�_^[�Ë�U���,�Pg3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�8�  3ۃ�;�u����SSSSS�0�J��������Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P�f�  ��;�t���u�E�SV�u���`������M�_^3�[�W����Ë�U���0�Pg3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�}�  3ۃ�;�u�d���SSSSS�8菜�������   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW诤  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[�]����Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3����o�6������Y���(r�_^Ë�Vh   h   3�V�v�  ����tVVVVV�ƙ����^Ë�U�������]�����]��E��u��M��m��]����]�����z3�@��3���h�������th��P�|���tj �������U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]Ã%�� Ë�U��3�9Ej ��h   P��������u]�3�@�|�]Ã=|�uWS3�9d�W�=P�~3V�5h���h �  j �v�����6j �5���׃�C;d�|�^�5h�j �5����_[�5������%�� Ë�VW3�����<�pu��p�8h�  �0���1�  YY��tF��$|�3�@_^Ã$�p 3����S�$�V�pW�>��t�~tW��W�~����& Y����0q|ܾp_���t	�~uP�Ӄ���0q|�^[Ë�U��E�4�p�,�]�jh�N�  3�G�}�3�9��u�s;  j��9  h�   �=  YY�u�4�p9t���nj袺��Y��;�u�#����    3��Qj
�Y   Y�]�9u,h�  W�(�  YY��uW謗��Y������    �]���>�W著��Y�E������	   �E��F  �j
�(���YË�U��EV�4�p�> uP�"���Y��uj�<  Y�6�(�^]Ë�U��d��h�k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �H�����   �x��5��h @  ��H� �  SQ�֋x��H��   ���	P�H��@�x�����    �H��@�HC�H��H�yC u	�`��H��x�ueSj �p�֡H��pj �5���P��d��H�k��h�+ȍL�Q�HQP�ˋ���E���d�;H�v�m�h��p��E�H��=x�[_^�át�V�5d�W3�;�u4��k�P�5h�W�5�����;�u3��x�t��5d��h�k�5h�h�A  j�5���`��F;�t�jh    h   W����F;�u�vW�5���P�뛃N��>�~�d��F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�����u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U����d��Mk�h�������M���SI�� VW}�����M���������3���U��p�����S�;#U�#��u
���];�r�;�u�h���S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1�h��	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t�p��C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;H�u�M�;x�u�%H� �M���B_^[��h�d�5    �D$�l$�l$+�SVW�Pg1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q���������������̋�U���S�]V�s35PgW��E� �E�   �{���t�N�38��~���N�F�38��~���E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���p�  �E���|@G�E��؃��u΀}� t$����t�N�38�P~���N�V�3:�@~���E�_^[��]��E�    �ɋM�9csm�u)�=,� t h,�胗  ����t�UjR�,����M��  �E9XthPgW�Ӌ���  �E�M��H����t�N�38�}���N�V�3:�}���E��H��詍  �����9S�R���hPgW�����  �����0qá`�Vj^��u�   �;�}�ƣ`�jP�Y���YY�@���ujV�5`��@���YY�@���ujX^�3ҹ0q��@���� �����s|�j�^3ҹ@qW������@�����������t;�t��u�1�� B���q|�_3�^�詏���=�� t��  �5@�貉��YË�U��V�u�0q;�r"���sw��+�����Q�����N �  Y�
�� V�(�^]Ë�U��E��}��P������E�H �  Y]ËE�� P�(�]Ë�U��E�0q;�r=�sw�`���+�����P�����Y]Ã� P�,�]Ë�U��M���E}�`�����Q����Y]Ã� P�,�]Ë�U��V�uW3�;�u����WWWWW�    �+�������   �F����   �@��   �t�� �F��   ���F�  u	V�  Y��F��v�vV�W  YP���  ���F;���   �����   �F�uOV�-  Y���t.V�!  Y���t"V�  ��V�<�@��  ��Y��Y���s�@$�<�u�N    �~   u�F�t�   u�F   ��N�A���������	F�~���_^]�jThO� ���3��}��E�P����E�����j@j ^V�y���YY;��  �@��5(���   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@�@���   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M���@���(� ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=(�|���=(��e� ��~m�E����tV���tQ��tK�uQ�����t<�u���������4�@��E� ���Fh�  �FP蟑  YY����   �F�E�C�E�9}�|�3ۋ���5@�����t���t�N��r�F���uj�X�
��H������P��������tC��t?W�����t4�>%�   ��u�N@�	��u�Nh�  �FP�	�  YY��t7�F�
�N@�����C���g����5(����3��3�@Ëe��E������������Ë�VW�@��>��t1��   �� t
�GP�$����@   ;�r��6�����& Y����@�|�_^Ë�U��EV3�;�u�8���VVVVV�    �_����������@^]Ë�U��QV�uV�����E�FY��u������ 	   �N ����/  �@t������ "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,������� ;�t�������@;�u�u�`�  Y��uV��   Y�F  W��   �F�>�H��N+�I;��N~WP�u�  ���E��M�� �F����y�M���t���t�����������@����s�@ tjSSQ���  #����t%�F�M��3�GW�EP�u�  ���E�9}�t	�N �����E%�   _[^�Ë�U���L�h   ����Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U���  ��  �Pg3ŉE��EV3���4�����8�����0���9uu3���  ;�u'�:����0� ���VVVVV�    �G���������  SW�}�����4�@������ǊX$�����(�����'�����t��u0�M����u&�����3��0����VVVVV�    �܁�����C  �@ tjj j �u�ʖ  ���u�]�  Y����  ��D���  ������@l3�9H�������P��4�� ���������`  3�9� ���t���P  �����4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P��  Y��t:��4���+�M3�@;���  j��@���SP覙  �������  C��D����jS��@���P肙  �������  3�PPj�M�Qj��@���QP�����C��D����h������\  j ��<���PV�E�P��(���� �4������)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4�������  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@���菖  Yf;�@����h  ��8����� ��� t)jXP��@����b�  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4������B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4������b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �h���;���   j ��,���P��+�P��5����P��(���� �4�����t�,���;����L���@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0�����t��,�����@��� ��8�����L���@�����8��� ul��@��� t-j^9�@���u����� 	   �����0�?��@�������Y�1��(�����D@t��4����8u3��$�h����    �p����  ������8���+�0���_[�M�3�^��n����jh(O�l����E���u�4����  ����� 	   ����   3�;�|;(�r!�����8������ 	   WWWWW�{�����ɋ�����@���������L1��t�P�m�  Y�}���D0t�u�u�u�.������E������� 	   �����8�M���E������	   �E��������u跕  Y�jhHO�����E���u�E���� 	   ����   3�;�|;(�r�$���� 	   SSSSS�Kz�����Ћ����<�@���������L��t�P蠔  Y�]���Dt1�u��  YP�����u�L��E���]�9]�t������M������ 	   �M���E������	   �E�������u�֔  YË�U��V�u�F��t�t�v�z���f����3�Y��F�F^]Ë�U��   ��~  �Pg3ŉE�SV�uWV�������3�9FY������}�FjPPS�Ў  ������������������|��s
������  ������@���������� ��ÊH$����F  ������u�F�������+�ʋǋ��  ��V��+��V���������Z  �������  3�9P0�  �����9Vu�������������<  R�p,�p(���������  ��������� Ã���;p(�0���;x,�'���j ������Qh   ������Q�0���������j ������������������融  ����������������������������;��������������t7������K;�s+���u�J�;�s�H�9
u�������`w�@��uЍ�����+�3����L  �@�t�V��:
u������B;�r������������u�������  ��x������    �$����F��   �V��u!�������   +N��@�����   jj j ������蛌  ��;�����u$;�����u�F�8��8
uG@;�r��F    �Yj �������������������S�  �����������������   ;�w�N��t
����   t�~������� �DtG������u��)����������� ������uѭ����������3������������M�_^3�[�i����jhhO�2����u�����Y�e� �u����Y�E��U��E������   �E��U��D�����u�4���YË�U��V�uV��  Y���u����� 	   ����MW�uj �uP��������u�L��3���tP����Y����������@������D0� ���_^]�jh�O�s����E���u�;����  � ���� 	   ����   3�;�|;(�r!�����8������ 	   WWWWW�u�����ɋ�����@���������L1��t�P�t�  Y�}���D0t�u�u�u��������E������� 	   �����8�M���E������	   �E��������u辏  YË�U���SW�}3�;�u �M���SSSSS�    �tt��������f  W�����9_Y�E�}�_jSP�������;ÉE�|ӋW��  u+G�.  ��OV��+�u���tA�U��u�����@������D2�t��;�s���:
u�E�3�B;�r�9]�u�E���   ��x������    �   �G��   �W;�u�]��   �]��u�+��������@��E����D0�tyjj �u�������;E�u �G�M��	�8
u�E@;�r��G    �@j �u��u����������}����:�   9Ew�O��t��   t�G�E��D0t�E�E)E��E�M��^_[�Ë�U��V�u�FW��ty�}��t
��t��uh���F��uV�I���EYU3�V�@w���FY��y����F��t�t�   u�F   W�u�uV����YP��  #����t3���9����    ���_^]�jh�O�^����u�!���Y�e� �u�u�u�u�:������E��E������	   �E��k�����u�[���YË�U��V�uWV��  Y���tP�@���u	���   u��u�@Dtj��  j���ً  YY;�tV�͋  YP� ���u
�L����3�V�)�  ������@�����Y�D0 ��tW�s���Y����3�_^]�jh�O�s����E���u�;����  � ���� 	   ����   3�;�|;(�r!�����8������ 	   WWWWW�q�����ɋ�����@���������L1��t�P�t�  Y�}���D0t�u�����Y�E������� 	   �M���E������	   �E�������u�͋  YË�U��9EuF�jP;Mu+����YY���u3�]ËE�    �6�u�7�~������Q��������tՉ�&3�@]Ë�U���EP�`������EYu��߃�]��Jx	�
�A�
�R�����YË�U��}�t]�-s��]Ë�U��S�U�������؃��t��P����Y��u��[]Ë�U����  �Pg3ŉE��M�EV3�W�}�������|�����d�����T���ǅ$���^  ��0����������x���;�u �K���VVVVV�    �ro��������5  ;�t��@@SuzP�����Y��s���t���t�ȃ��������@�����A$u&���t���t�ȃ������@�����@$�t �����VVVVV�    ��n��������  �u�������b���ƅc��� ��t�����<������k  ��d�����P�ȍ��Y��t0��t���VV��t�������YP�k���YYG�P蝍��Y��u��  �<%�1  8G�  3���@���ƅ/��� ��X�����L�����l���ƅa��� ƅ`��� ƅj��� ƅS��� ƅb��� ƅs��� ƅk�����(���G���P����Y��t��l�����L���k�
�DЉ�l�����   ��N��   ��   ��*tp��F��   ��It��Lut��k����   �O��6u�G�84u��(�������4�����8����m��3u�G�82u���\��dtW��itR��otM��xtH��Xu�A��j����9��ht(��lt��wt��S����"�G�8lt���k�����s������k�����s�����S��� �������j��� ��H���u������0�������������3�2ۉ�D���8�s���u�<Stƅs����<Cuƅs������ ��\�����ntJ��ct��{t��d�����t����}���Y���d�����t����@�����x��������  ��D�����H�����L�����t��l��� ��  ��\�����o�r  �  ��c�
  jdZ;���  �z  ��g~E��it!��n�g  ��j��� ��t����f
  �
  ��\�����x���-�4  ƅ`����1  3ۃ�x���-u��T���� -C�	��x���+u��l�����d�����t����^�����x�����L��� u��l������x����k��l�����l�����tf��x�����T�����X������0���P��|���PCS��T�����$�������������
  ��d�����t����������x�����P����Y��u���������   � � ��a���:�x�����   ��l�����l�������   ��d�����t���������T�����x�����a������0���P��|���PCS��T�����$��������������	  ��x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$����{���������	  ��d�����t����������x�����P����Y��u���X��� �_  ��x���et��x���E�I  ��l�����l������5  ��T����e��0���P��|���PCS��T�����$��������������  ��d�����t����D�����x�����-u,��T����-��0���P��|���PCS����������  �	��x���+u/��l�����l�����u!�l������d�����t����������x�����x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$������������  ��d�����t����j�����x�����P誆��Y��u���d�����t�����x����U�����X��� YY��  ��j��� ��  ��T�����<��������QP��D���� ��k���HP�5�o�&���Y�Ѓ��  ��u��l���ǅL���   ��s��� ~ƅb�����d�����t���W��x�����@�������YY��L��� t��l�����l������3  ��t������x�����x�������  ��\���ctN��\���su��	|	����  �� u2��\���{��  ��a���3ҋȃ�B������L�3˅���  ��j��� ��  ��b��� �~  �� �����P�#k  Y��t��t������������!��������P�����ǅ���?   ���   �� ���P�����P�~  f�������f�FF�  ��p��  �������HH�{  ���������t3�;�x�����  ��c�����j��� �  �����������  ��s��� ~ƅb���G�?^��u
�wƅa����j �E�j P�V]�����>]u	�]F�E� �f��/����^F<-uB��t>���]t7F:�s�����:�w"*������Ћσ��ǳ�����D�GJu�2���ȊЋ��������D��<]u����  ��H�����D���������x���+u'��l���u��t����d�����t����C�����x���j0^9�x����x  ��d�����t���������x���<xtX<XtT��\���xǅX���   t"��L��� t
��l���u��ǅ\���o   �$  ��d�����t���P�����YY��x����  ��d�����t���������L��� ��x���t��l�����l���}��ǅ\���x   ��   �F��D����������@���������t���WP�j���YY9�@�����  ��j��� �  ��<�����\���c��  ��b��� t��D���3�f���  ��D����  ��  ƅk�����x���-u	ƅ`����	��x���+u'��l���u��t����d�����t���������x�����(��� �J  ���  ��\���xte��\���pt\��x���P�с��Y����   ��\���ou"��x���8��   ��4�����8��������Rj j
��8�����4�����^�������7��x���P�����Y��tr��4�����8�����x������������Y��x�����x�����X�����Й����L��� ��4�����8���t��l���t5��d�����t���������x���������d�����t�����x�������YY��`��� ��@�����   ��4�����8����؃� �ى�4�����8�����   ��@�������   ��\���xt;��\���pt2��x���P聀��Y����   ��\���ou��x���8}n���,k�
�'��x���P�Ӏ��Y��tR��x����������Y��x�����X�����L��� ��x����|�t��l���t5��d�����t���������x����X�����d�����t�����x�������YY��`��� t�߃�\���Fu��X��� ��X��� �  ��j��� u8��<�����D�����(��� t��4������8����F���k��� t�>�f�>��H�����c���G��H����`<%u
�G�8%u����t�������������G��x�����H���;�ul��P�e  Y��t!��t�����������G��H���;�uG��t�����x����u�?%uD��H����xnu8������	����*��d�����x�������YY�VS��VP����VS�y�������0���u��T����a��Y��x����u*��<�����u8�c���u�������� t%������ap������� t
������`p���<���[�M�_3�^�S���Ë�U���VW�u�M��
T���E�u3�;�t�0;�u,�����WWWWW�    ��_�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�4*  �M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&� ����E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9luh`n�P������]Ë�U��QQS�]VW3�3��}�;��st	G�}���r���w  j�|  Y���4  j�p|  Y��u�=`�  ���   �A  h��  S�P�W� T������tVVVVV�\����h  �i�Vj �m� �����u&h�h�  V�S������t3�PPPPP��[����V�`���@Y��<v8V�S�����;�j�d�h�+�QP�/<  ����t3�VVVVV�[�����3�h�SW�E;  ����tVVVVV�k[�����E��4��sSW� ;  ����tVVVVV�F[����h  h`W��y  ���2j������;�t$���tj �E�P�4��s�6螀��YP�6S���_^[��j�{  Y��tj��z  Y��u�=`uh�   �)���h�   ����YYË�U���   �Pg3ŉE��ESV�u3ۃ}W��t�����l�����   Sh�   ��|�����Q�u��x����uP�:|  ����;�uj�L���z��   SSS�u�u��t����|  ����p���;�t_3�FVP��~����YY;�tMS��p�����x���W�u�u��t�����{  ����;�tjV�~��YY��l����;�u!9�x���tW�z[��Y����M�_^3�[�bN���ÍN�QWVP�>:  ����tSSSSS�Y����9�x���tW�9[��Y3��9]u�Sj�d�W�u�uP��y  ����t�����P�x��Y��tɊ�
���,0GG��l��|�뱋�U��E�l�]Ë�U��W��  W���u�x����  ��`�  w��t�_]Ë�U��������u�L����5�t����h�   �Ѓ�]Ë�U��h��x���th�P�|���t�u��]Ë�U���u�����Y�u����j�����Y�j�����YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=H� thH��@f  Y��t
�u�H�Y����h��hx�����YY��uBh���p���\��$t��c����=$� Yth$���e  Y��tj jj �$�3�]�jh�O�����j�����Y�e� 3�C9����   ����E����} ��   �5�蛠��Y���}؅�tx�5�膠��Y���u܉}�u����u�;�rW�b���9t�;�rJ�6�\������L�������5��F������5��9�����9}�u9E�t�}�}؉E����u܋}��h������_���Yh������O���Y�E������   �} u(���j����Y�u�����3�C�} tj�����Y�����Ë�U��j j�u�������]�jj j ������Ë�V胟����V�
  V�`c  V�@V��V�
���V�Sx  V�e(  V��  V�n���h���՞����$��t^Ã= � u胮��V�5TW3���u����   <=tGV�{��Y�t���u�jGW�z����YY�=����tˋ5TS�BV�T{����C�>=Yt1jS�Uz��YY���tNVSP�uM������t3�PPPPP�U�������> u��5T�W���%T �' ��   3�Y[_^��5����V���%�� ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�Ww  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�rv  Y��t��M�E�F��M��E���Ov  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9 �u�����h  ���VS����������5��;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�w����Y;�t)�U��E�P�WV�}�������E���H�t��5x�3�����_^[�Ë�U�조���SV�5��W3�3�;�u.�֋�;�t���   �#�L���xu
jX�����������   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5h�SSS+�S��@PWSS�E��։E�;�t/P�v��Y�E�;�t!SS�u�P�u�WSS�օ�u�u���S��Y�]��]�W������\��t;�u������;��r���8t
@8u�@8u�+�@P�E��Ev����Y;�uV����E����u�VW��e����V�����_^[�Ë�V��%��%W��;�s���t�Ѓ�;�r�_^Ë�V��%��%W��;�s���t�Ѓ�;�r�_^�Ë�U��QQV�U��������F  �V\��tW�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ��t�=�t���;�}$k��~\�d9 �=�t��tB߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]Ë�U����Pg�e� �e� SW�N�@��  ��;�t��t	�УTg�`V�E�P���u�3u�� �3��X�3����3��E�P����E�3E�3�;�u�O�@����u������5Pg�։5Tg^_[�Ë�U���(3�S�]V�uW�}�E��E��E��E��E��E��E��E�9��t�5��8���Y��!�M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E�$��M��]�Q��]���]���Y����  �m���� "   �  �E� ��M��]�Q��E�   �]���]���Y�j  �E�   �E� ��E���]���]���"  �M��E��r����E��׉M��E��Z����E�$놃�tNIt?It0It ��t����   �E���E���E�$����E�$�x����E�   ��������   �E�   �E����������������   �$����E���E���E� ��E����E����E���y����E���m����E����E����E����M����]���]�M��]�Q�E�   ��Y��u�ե��� !   �E��_^[�������������%�����1�:�C��%� �=�����3�Ë�U��QQSV���  V�5�t�vw  �EYY�M�ظ�  #�QQ�$f;�uU�v  YY��~-��~��u#�ESQQ�$j�t  ���rVS�*w  �EYY�d�ES�h����\$�E�$jj�?�u  �]��EY�]�Y����DzVS��v  �E�YY�"�� u��E�S���\$�E�$jj�t  ��^[�Ë�U��E���]Ë�U���5�������Y��t�u��Y��t3�@]�3�]Ë�U��� S3�9]u �\���SSSSS�    �L��������   �MV�u;�t!;�u�-���SSSSS�    �TL��������S�����E�;�w�M�W�u�E��u�E�B   �u�u�P�u��w  ����;�t�M�x�E����E�PS����YY��_^[�Ë�U���uj �u�u�u�5�����]�jhP�ӿ��3��]3�;���;�u耣���    WWWWW�K��������S�=|�u8j蟴��Y�}�S�ȴ��Y�E�;�t�s���	�u���u��E������%   9}�uSW�5��������蓿���3��]�u�j�m���Y�����U���0���S�ٽ\�����=px t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=px t�#  ��8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����,  �   [�À�8�����=D uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �H�����������8����s4�X�,ǅr���   �@�����������0����v�PVW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�:�  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����D   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Àzuf��\���������?�f�?f��^���٭^�����t�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����t�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����t���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-�t��p��� ƅp���
��
�t����������l$�l$�D$���   5   �   t��������t u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t� u��� u���l$����u���u���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r �������u�|$�l$�ɛ�l$������l$��Ã�,��?�$�Nu����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  ������u �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����<u�Ƀ�u�\$0�|$(���l$�-Du�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�,u�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���$u�|$�$u�<$� �|$$�D$$   �D$(�l$(���$u�<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  ������u �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����<u�Ƀ�u�\$0�|$(���l$�-Du�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8�,u�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w���$u�|$�$u�<$� �|$$�D$$   �D$(�l$(���$u�<$�l$$�Q�����0Z�����0Z�������@���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�p  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��`�   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��������������|�����   s�����������������t�����   v���떋�U����Pg3ŉE�j�E�Ph  �u�E� ����u����
�E�P�D��Y�M�3��*���Ë�U���4�Pg3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5t��M�QP�֋l���t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u��[����YF;�~[�����wS�D6=   w/蔎����;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�~H��Y;�t	� ��  ���E���}�9}�t؍6PW�u��<-����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�h���t`�]��[�h�9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�;Y��YY�E�;�t+WWVPV�u�W�u��;�u�u��6��Y�}���}��t�MЉ�u��Y)��Y�E��e�_^[�M�3���(���Ë�U���S�u�M��O)���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P��8  YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP��  �� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U��QQ�Pg3ŉE����SV3�W��;�u:�E�P3�FVh �V����t�5���4�L���xu
jX�����������   ;���   ����   �]�9]u��@�E�5l�3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w������;�t� ��  �P�	F��Y;�t	� ��  ���؅�ti�?Pj S��*����WS�u�uj�u�օ�t�uPS�u���E�S�^'���E�Y�u3�9]u��@�E9]u��@�E�u�����Y���u3��G;EtSS�MQ�uP�u��������;�t܉u�u�u�u�u�u����;�tV�3��Y�Ǎe�_^[�M�3��s&���Ë�U����u�M���&���u$�M��u �u�u�u�u�u�������}� t�M��ap���jh(P详���M3�;�v.j�X3���;E�@u�T����    WWWWW�{2����3���   �M��u;�u3�F3ۉ]���wi�=|�uK������u�E;l�w7j�C���Y�}��u�I���Y�E��E������_   �]�;�t�uWS�%)����;�uaVj�5���`���;�uL9=��t3V����Y���r����E;��P����    �E���3��uj����Y�;�u�E;�t�    �������jhHP葥���]��u�u�C��Y��  �u��uS��1��Y�  �=|���  3��}�����  j�P���Y�}�S�y���Y�E�;���   ;5l�wIVSP�[�������t�]��5V�*���Y�E�;�t'�C�H;�r��PS�u���C��S�)����E�SP�O�����9}�uH;�u3�F�u������uVW�5���`��E�;�t �C�H;�r��PS�u��C��S�u��������E������.   �}� u1��uF������uVSj �5���������u�]j聘��YË}����   9=��t,V�`���Y�����������9}�ul���L�P薇��Y��_����   �Ƈ��9}�th�    �q��uFVSj �5���������uV9��t4V�����Y��t���v�V�����Y�z����    3�������g����|�����u�Y������L�P�	����Y���ҋ�U��MS3�;�v(j�3�X��;Es�$���SSSSS�    �K/����3��A�MVW��9]t�u�W���Y��V�u������YY��t;�s+�Vj �S�)&������_^[]Ë�U��E�Ĉ�Ȉ�̈�Ј]Ë�U��E��tV9Pt��k�u��;�r�k�M^;�s9Pt3�]��5̈�v��Y�j hhP虢��3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�:x�����}؅�u����a  �Ĉ�Ĉ�`�w\���]���������Z�Ã�t<��t+Ht�����    3�PPPPP�.����뮾̈�̈��Ȉ�Ȉ�
�Ј�Ј�E�   P��u���E�Y3��}���   9E�uj����9E�tP�Ŗ��Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.��t�M܋�t��t�9M�}�M�k��W\�D�E����Eu����E������   ��u�wdS�U�Y��]�}؃}� tj �S���Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3��;���Ë�U����HB�PD�M��U���u����Ãe� SW�E��FPj1Q3�C�E�SP��������FPj2�u��E�SP������FPj3�u��E�SP������FPj4�u��E�SP������P��FPj5�u��E�SP�u�����FPj6�u��E�SP�`���Vj7�u���E�SP�N�����F Pj*�u��E�SP�9�����P��F$Pj+�u��E�SP�!�����F(Pj,�u��E�SP������F,Pj-�u��E�SP�������F0Pj.�u��E�SP�������P��F4Pj/�u��E�SP�������FPj0�u��E�SP������F8PjD�u��E�SP������F<PjE�u��E�SP������P��F@PjF�u��E�SP�s�����FDPjG�u��E�SP�^�����FHPjH�u��E�SP�I�����FLPjI�u��E�SP�4�����P��FPPjJ�u��E�SP������FTPjK�u��E�SP������FXPjL�u��E�SP�������F\PjM�u��E�SP�������P��F`PjN�u��E�SP�������FdPjO�u��E�SP������FhPj8�u��E�SP������FlPj9�u��E�SP������P��FpPj:�u��E�SP�n�����FtPj;�u��E�SP�Y�����FxPj<�u��E�SP�D�����F|Pj=�u��E�SP�/�����P����   Pj>�u��E�SP��������   Pj?�u��E�SP���������   Pj@�u�S�E�P���������   PjA�u��E�SP�������P����   PjB�u��E�SP��������   PjC�u��E�SP��������   Pj(�u��E�SP��������   Pj)�u��E�SP�i�����P����   Pj�u��E�SP�N�������   Pj �u��E�SP�6�������   Ph  �u��E�SP��������   Ph	  �]�S�E�j P�������P���_���   [�Ë�U��V�u����  �v�<)���v�4)���v�,)���v�$)���v�)���v�)���6�)���v �)���v$��(���v(��(���v,��(���v0��(���v4��(���v��(���v8��(���v<��(����@�v@�(���vD�(���vH�(���vL�(���vP�(���vT�(���vX�(���v\�(���v`�z(���vd�r(���vh�j(���vl�b(���vp�Z(���vt�R(���vx�J(���v|�B(����@���   �4(�����   �)(�����   �(�����   �(�����   �(�����   ��'�����   ��'�����   ��'�����   ��'�����   ��'�����   ��'����,^]Ë�U��SVW�}�  �Pvt@h�   j�J����YY��u3�@�E��������tV�+���V�z'��YY��ǆ�      �����   �;�t�   P���73�_^[]Ë�U��V�u��t5�;wtP�*'��Y�F;wtP�'��Y�v;5wtV�'��Y^]Ë�U���S�]V3�W�]�u�9su9su�u��u��Ew�:  j0j��I����YY�};�u3�@�w  ���   jYj��\I��3�Y�E�;�u�u�&��Y�щ09s��   j�5I��Y�E�;�u3�F�u�h&���u��`&��YY���  �0�u�{>VjW�E�jP������E�FPjW�E�jP�����	E�FPjW�E��E�jP������<E�tV����Y���뎋E�� ����0|��9��0�@�8 u��7��;u���~�����> u���w�E��w�H�w�u��H�E�3�A��E���t����   �5���tP�֋��   ��tP�օ�u���   �g%�����   �\%��YY�E����   �E����   �E���   3�_^[�Ë�U��V�u��t~�F;wtP�%��Y�F; wtP�%��Y�F;$wtP��$��Y�F;(wtP��$��Y�F;,wtP��$��Y�F ;0wtP��$��Y�v$;54wtV�$��Y^]Ë�U���SV�uW3��}��u��}�9~u9~u�}��}��w�6  j0j�mG����YY;�u3�@�u  j�G��Y�E�;�u	S�I$��Y���89~��  j��F��Y�E�;�uS�&$���u��$��Y�҉8�v8�CPjV�E�jP�������CPjV�E�jP������CPjV�E�jP�s�����CPjV�E�jP�_�����P��CPjV�E�jP�H�����C PjPV�E�jP�4�����C$PjQV�E�jP� �����C(PjV�E�j P������P��C)PjVj �E�P�������C*PjTV�E�j P�������C+PjUV�E�j P�������C,PjVV�E�j P������P��C-PjWV�E�j P������C.PjRV�E�j P������C/PjSV�E�j P�z�����<�t$S����S��"���u���"���u��"�����Q����C����0|��9��0�@�8 u��#��;u���~�����> u���jY�w���E�u�   ��	���I�K� �@�M��C3�@3��9}�t�M�����   ;�tP�����   ;�t#P����u���   �"�����   �"��YY�E����   �E����   ���   3�_^[��3�Ë�U��ES3�VW;�t�};�w�y��j^�0SSSSS�3!�������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u���x��j"Y����3�_^[]�����������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^�Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w�2x��j^�0SSSSS�Z ��������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x�����w��j"Y���낋�U��3�S3�@9]|FVW��t>�EÙ+��E���<��7�E�0�Y  YY��u
�M���9�}N�u��^;]~�_^3Ʌ���[��]Ë�U����Pg3ŉE�V���tS�> tNh�V�Zo��YY��t=h�V�Io��YY��uj�E�Pj�w����t/�u�V�,��Y�M�3�^�����j�E�Ph  �w����u3��׍E�h�P��n��YY��u����뻋�U��3�f�Mf;��t@@��r�3�@]�3�]Ë�V3��#��,aB<w������,A<w��������tЊ
��u׋�^�3��
B��A|��Z~��a��w@��Ë�U���|�Pg3ŉE�VW�}�h�����ׁƜ   ������jx�E�P�F���%���  PW����u!F@�2�E�P�v�eW  YY��uW����Y��t
�N�~�~�F���Ѓ��M�_3�^�T���� ��U���|�Pg3ŉE�Vjx�E�P�E%�  j   P������u3��.�U������9Et�} t�6W�������V����A��Y;�_t�3�@�M�3�^�����Ë�U���|�Pg3ŉE�SVW�}�g�����ׁƜ   �y�������jx�E�P�F���%���  PW�Ӆ�u�f 3�@�b  �E�P�v�PV  YY����   jx�E�P�F���%���  PW�Ӆ�t��E�P�6�V  YY��u�N  �~�R�FuO�F��t,P�E�P�6�5W  ����u�6�N�~��@��Y;Fu!�~��V��uW����Y��t	���V�~�N�   #�;���   jx�E�P�F���%���  PW�Ӆ������E�P�6�uU  Y3�Y��u/�N   �F9^t
   �F�G9^t;�6�]@��Y;Fu.j�9^u49^t/�E�P�6�)U  YY��uSW�������YY��t�N   9^u�~�F���Ѓ��M�_^3�[����� ��U���|�Pg3ŉE�VW�}��e�����ׁƜ   ������jx�E�P�F���%���  PW����u!F@�[�E�P�6�T  YY��u	9Fu0j��~ u0�~ t*�E�P�6�bT  YY��uPW���$���YY��t
�N�~�~�F���Ѓ��M�_3�^�M���� �6�6?���v�����@�F�#?��������f @�~ YY�FtjX���	���jh %�F���F�   t�   t�u�f ��6��>�������@Y�FtjX������jh�&�F���Fu�f Ë�U��SVW�kd���]���Ɯ   ��u�N  �   �C@�~����t�8 tWjh����������f ��tS�8 tN���t�8 t�������S����~ ��   Vj@h�	��������tb�?��t�? t�����P�����I�?��t0�? t+W��=������Y�j@h$�F���Fu�f ��F  ���F�F�~ ��   �˃����#ˋ��������}����   ����  ��   ����  ��   ��P�������   j�v� �����   �E��tf�Nf�f�Nf�Hf�x�]��tm�=��  f9u%h�j@S�G������t"3�PPPPP�[�����j@Sh  �v�ׅ�t,j@�C@Ph  �v�ׅ�tj
j��S�u�"T  ��3�@�3�_^[]Ë�U��VW�}�ǃ� ��  H��  H��  H�I  H��  �M�ESj Z�r  �0;1t|�0�+�t3ۅ��Í\�����i  �p�Y+�t3ۅ��Í\�����H  �p�Y+�t3ۅ��Í\�����'  �p�Y+�t3ۅ��Í\����3����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3����r  �p;qt~�p�Y+�t3ۅ��Í\�����I  �p	�Y	+�t3ۅ��Í\�����(  �p
�Y
+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����w  �p�Y+�t3ۅ��Í\����3����R  �p;qt~�Y�p+�t3ۅ��Í\�����)  �p�Y+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����x  �p�Y+�t3ۅ��Í\�����W  �p�Y+�t3ۅ��Í\����3����2  �p;qt~�p�Y+�t3ۅ��Í\�����	  �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\����3�����   �p;qtr�p�Y+�t3ۅ��Í\����u}�p�Y+�t3ۅ��Í\����u`�p�Y+�t3ۅ��Í\����uC�p�Y+�t3ۅ��Í\����3���u"��+�;�������σ���  �$�G@����  �P�;Q�tq���Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����3����v����P�;Q�t}���Q�+�t3҅��T�����N����p��Q�+�t3҅��T�����-����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����}����p��Q�+�t3҅��T����3����X����P�;Q�t}���Q�+�t3҅��T�����0����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T�����^����p��Q�+�t3҅��T����3����9����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�to���Q�+�t3҅��T���u6�p��Q�+�t3҅��T���u�p��Q�+�t3҅��T���t����@��I�+�t3Ʌ����L	����3���u3�[�S  �P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����n����p��Q�+�t3҅��T�����M����p��Q�+�t3҅��T�����,����p��Q�+�t3҅��T����3��������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����x����P�;Q�t}���Q�+�t3҅��T�����P����p��Q�+�t3҅��T�����/����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3����Z����P�;Q�t~�Q��p�+�t3҅��T�����1����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����`����p��Q�+�t3҅��T����3����;����I��@�+�� ���3Ʌ����L	���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����b����p��Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����l����P�;Q�t}���Q�+�t3҅��T�����D����p��Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����s����p��Q�+�t3҅��T����3����N����P�;Q�t~�Q��p�+�t3҅��T�����%����Q��p�+�t3҅��T���������Q��p�+�t3҅��T����������Q��p�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T����3����/���f�P�f;Q�������Q��p�+������3҅��T����  �����P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����i����P�;Q�t}���Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����p����p��Q�+�t3҅��T����3����K����P�;Q�t}���Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T�����r����p��Q�+�t3҅��T�����Q����p��Q�+�t3҅��T����3����,����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T�����3����p��Q�+�t3҅��T����3��������p��Q�+������3҅��T���������������M�u��+�t3҅��T�����   �A�V+�t3҅��T�����   �A�V+�t3҅��T�����   �A�N+���   3Ʌ����L	����   �M�u��+�t3҅��T���uh�A�V+�t3҅��T���uK�A�N랋M�u��+�t3҅��T���u �A�N�p����E�M� �	�_���3�_^]��2�6�:?k2K6W:x>�1�5�9�=L1,589Y=�0�4�8�<.048;<�/3�7�;/�2�6;���������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U������SV�uW3��E��}�}��}��FFf�> t����at8��rt+��wt��X��WWWWW�    �����3��S  �  �3ۃM��	�	  �M�3�AFF�f;���  � @  ;��   ����S��   ��   �� ��   ��tVHtG��t1��
t!���u���9}���   �E�   ����   �ˀ   �   ��@��   ��@�   �E�   �   ����   �E����������   �E��}9}�ur�E�   �� �l��TtX��tCHt/��t��������� �  uC��E9}�u:�e������E�   �09}�u%	U��E�   ��� �  u�� �  ��   ��t3���FF�f;������9}���   �FFf�> t�jVh��>E  �����`���j ��X�FFf9t�f�>=�G���FFf9t�jh�V�`D  ����u��
��   �Djh�V�AD  ����u����   �%jh�V�"D  �������������   �FFf�> t�f9>�����h�  �u�ES�uP��B  ����������E�L��M��H�M�x�8�x�x�H_^[��jh�P�r��3�3��}�j�g��Y�]�3��u�;5`���   �@���9t[� �@��uH� �  uA�F���w�FP�f��Y����   �@��4�V�]u��YY�@����@�tPV�u��YYF둋��}��h��j8�Y!��Y�@���@��9tIh�  � �� P��	  YY���@�u�4�g���Y�@������ P�(��@��<�}�_;�t�g �  �_�_��_�O��E������   ����q��Ë}�j�e��Y�SVW�T$�D$�L$URPQQh�Ed�5    �Pg3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�R  �   �C�d  �d�    ��_^[ËL$�A   �   t3�D$�H3��P���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�  3�3�3�3�3���U��SVWj j h3FQ�i  _^[]�U�l$RQ�t$������]� ��U����u�M������E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U��3�@�} u3�]�U��SVWUj j h�F�u�i  ]_^[��]ËL$�A   �   t2�D$�H�3�����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�Fd�5    �Pg3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�Fu�Q�R9Qu�   �SQ�Pw�SQ�Pw�L$�K�C�kUQPXY]Y[� ����������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �������U��W�}3�������ك��E���8t3�����_�Ë�U���SV�u�M������]�   ;�sT�M胹�   ~�E�PjS�����M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�h���YY��t�Ej�E��]��E� Y��FQ��� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�����$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=l u�E�H���w�� ]�j �u�����YY]Ë�U���(�Pg3ŉE�SV�uW�u�}�M�������E�P3�SSSSW�E�P�E�P�I  �E�E�VP�?  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[������Ë�U���(�Pg3ŉE�SV�uW�u�}�M�� ����E�P3�SSSSW�E�P�E�P��H  �E�E�VP�C  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[� ����Ë�U��MSV�u3�W�y;�u�PO��j^�0SSSSS�x��������   9]v݋U;ӈ~���3�@9Ew�O��j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�f��@PWV������3�_^[]Ë�U��Q�M�ASVW������  #�% �  �߉E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��E��<  �U����������U��E�����P������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0�Pg3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f���M  �uЉC�E։�EԉC�E�P�uV�w�����$��t3�PPPPP�������M�_�s^��3�[�����������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�c���YË�U��E�M%����#�V������t1W�}3�;�tVV�V  YY��L��j_VVVVV�8�E�������_��uP�u��t	�bV  ���YV  YY3�^]Ë�U��E��]�jh�P�	h���e� �u�u�$��E��/�E� � �E�3�=  �����Ëe�}�  �uj����e� �E������E���g���������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h�Ph�d�    P��SVW�Pg1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh�P�Of��3ۉ]�j�L[��Y�]�j_�}�;=`�}W�����@��9tD� �@�tP����Y���t�E��|(�@���� P�$��@��4�a���Y�@��G��E������	   �E��f���j��Y��YË�U����UV�uj�X�E�U�;�u�pI���  �UI��� 	   ����  S3�;�|;5(�r'�FI����,I��SSSSS� 	   �S���������Q  ����W�<�@������ƊH��u� I�����H��� 	   �j�����wP�]�;��  ����  9]t7�@$����E���HjYtHu���Шt����U�E�E��   ���Шu!�H����zH���    SSSSS�������4����M;�r�E�u����Y�E�;�u�BH���    �JH���    ����h  jSS�u�^  ��D(�E���T,���AHtt�I��
tl9]tg��@�M�E�   �D
8]�tN��L%��
tC9]t>��@�M�}��E�   �D%
u$��L&��
t9]t��@�M�E�   �D&
S�M�Q�uP��4������{  �M�;��p  ;M�g  �M��D� ���  �}��  ;�t�M�9
u��� ��]�E�É]�E�;���   �M�<��   <t�CA�M�   �E�H;�s�A�8
u
AA�M�
�u�E�m�Ej �E�Pj�E�P��4�����u
�L���uE�}� t?��DHt�}�
t����M��L�%;]�u�}�
t�jj�j��u�  ���}�
t�C�E�9E�G������D� @u����C��+E�}��E���   ����   K���xC�   3�@�����;]�rK�@��`w t�����`w��u��E��� *   �zA;�u��@���AHt$C���Q|	���T%C��u	���T&C+���ؙjRP�u��  ���E�+]���P�uS�u�j h��  �l��E���u4�L�P�E��Y�M���E�;EtP����Y�E�����  �E��  �E��3�;�����E��L0��;�t�M�f�9
u��� ��]�E�É]�E�;���   �E�f����   f��tf�CC@@�E�   �M����;�s�Hf�9
u���Ej
�   �M�   �Ej �E�Pj�E�P��4�����u
�L���u[�}� tU��DHt(f�}�
t�jXf���M��L��M��L%��D&
�*;]�uf�}�
t�jj�j��u�|  ��f�}�
tjXf�CC�E�9E�������t�@u��f� f�CC+]�]������L�j^;�u��C��� 	   ��C���0�i�����m�Y����]��\���3�_[^��jhQ��_���E���u�C���  �C��� 	   ����   3�;�|;(�r!�C���0�sC��� 	   VVVVV�������ɋ�����@���������L9��t�����;M�Au�?C���0�%C���    �P��  Y�u���D8t�u�u�u�~������E����B��� 	   ��B���0�M���E������	   �E��M_����u�  YË�U��QQ�EV�u�E��EWV�E���  ���Y;�u�B��� 	   �ǋ��J�u�M�Q�u�P����E�;�u�L���t	P�B��Y�ϋ�����@������D0� ��E��U�_^��jh(Q�l^������u܉u��E���u�+B���  �B��� 	   �Ƌ���   3�;�|;(�r!�B���8��A��� 	   WWWWW�������ȋ�����@���������L1��u&��A���8�A��� 	   WWWWW�������������[P�=  Y�}���D0t�u�u�u�u�������E܉U���XA��� 	   �`A���8�M���M���E������   �E܋U��]����u�z  YË�U��E���u�A��� 	   3�]�V3�;�|;(�r��@��VVVVV� 	   ������3���ȃ�����@����D��@^]Ë�U����Pg3ŉE�V3�95`xtO�=�z�u�N  ��z���u���  �pV�M�Qj�MQP�0���ug�=`xu��L���xuω5`xVVj�E�Pj�EPV�,�P�h���z���t�V�U�RP�E�PQ�(���t�f�E�M�3�^�������`x   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M�������E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�l����E�u�M;��   r 8^t���   8]��e����M��ap��Y����"?��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�l����:���뺋�U��j �u�u�u�������]Ë�U��EVW��|Y;(�sQ���������<�@�����<�u5�=`S�]u�� tHtHuSj��Sj��Sj��4���3�[��[>��� 	   �c>���  ���_^]Ë�U��MS3�;�VW|[;(�sS������<�@��������@t5�8�t0�=`u+�tItIuSj��Sj��Sj��4����3����=��� 	   ��=������_^[]Ë�U��E���u��=���  �=��� 	   ���]�V3�;�|";(�s�ȃ�����@�����@u$�=���0�f=��VVVVV� 	   ����������� ^]�jhHQ�{Y���}����������4�@��E�   3�9^u6j
�XN��Y�]�9^uh�  �FP�#���YY��u�]��F�E������0   9]�t����������@��D8P�(��E��;Y���3ۋ}j
�M��YË�U��E�ȃ�����@����DP�,�]�jhhQ�X���M��3��}�j��L��Y��u����b  j�M��Y�}��}؃�@�<  �4�@�����   �u���@�   ;���   �Fu\�~ u9j
�PM��Y3�C�]��~ uh�  �FP����YY��u�]���F�e� �(   �}� u�^S�(��FtS�,���@낋}؋u�j
�L��YÃ}� u��F��+4�@���������u�}��uyG�+���j@j �(��YY�E���ta��@���(� ���   ;�s�@ ���@
�` ��@�E������}�����σ�����@��DW�����Y��u�M���E������	   �E��uW���j�WK��Y���������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U���SVW�d*���e� �= � ����   ht�8������*  �5|�hhW�օ��  P�)���$XW� ���P�)���$DW�$���P�)���$(W�(���P�o)��Y�0���thW��P�W)��Y�,��,�;�tO90�tGP�)���50����)��YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9�$�;�t0P�e)��Y��t%�ЉE���t�(�;�tP�H)��Y��t�u��ЉE��5 ��0)��Y��t�u�u�u�u����3�_^[�Ë�U��MV3�;�|��~��u�\�(�\�\��8��VVVVV�    ����������^]Ë�U����u�M������u�u�u�u�<��}� t�M��ap��Ë�U��QQ�Pg3ŉE��4�S�<�VW3�3�G;�u,VVWV�Ӆ�t�=4��/�L���xu
jX�4���4�����   ;���   ;�u#9uu�E� �@�EVV�u�u�ӋȉM�;�u3��   ~Ej�3�X���r9�D	=   w�8����;�t����  ���P����Y;�t	� ��  �����3�;�t��u�W�u�u�Ӆ�t VV9uuVV��u�uj�WV�u�h���W�Y���Y����u�u�u�u���e�_^[�M�3�������Ë�U����u�M��=����u�E��u�u�u�uP�������}� t�M��ap��Ë�U��E�8�]Ë�U����u�M�������E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u�H��M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�}  Y����  �t�Etj�c  Y����v  ����   �E��   j�A  �EY�   #�tT=   t7=   t;�ub��M����py��{L�H��M�����{,�py�2��M�����z�py���M�����z�`y��`y��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�x  �M��]�� �����������}�E���@��S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}�n1��� "   ]��a1��� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���xx;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P蔷������uV�,���Y�E�^�Ë�|x�h��  �u(�  �u�����E ���Ë�U��=px u(�u�E���\$���\$�E�$�uj�/�����$]��J0��h��  �u� !   �J  �EYY]Ë�S��QQ�����U�k�l$���   �Pg3ŉE��s �CP�s��������u"�e���CP�CP�s�C �sP�E�P�I������s�p������=px u+��t'�s �C���\$���\$�C�$�sP�r�����$�P�����$��  �s �  �CYY�M�3�� �����]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj���  f;�u�E�� u9Utj��3�]Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������"Q���EQQ�$����������  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�-�y�]���t����-�y�]�������t
�-�y�]����t	�������؛�� t���]����jh�Q�I��3�9��tV�E@tH9�yt@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�y �e��U�E�������e��U�~I����A@t�y t$�Ix��������QP�P��YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u�l,���8*u�ϰ?�d����} �^[]Ë�U���x  �Pg3ŉE�S�]V�u3�W�}�u������������������������������������������������������������������u5��+���    3�PPPPP�	����������� t
�������`p������
  �F@u^V�\O��Y��s���t���t�ȃ��������@�����A$u����t���t�ȃ������@�����@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw�������3��3�3����j��Y������;���	  �$�ny��������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�����������Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u��y������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P�d6  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  ��y������P�/���Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7����������3  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V�����������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5�o�>��Y�Ћ���������   t 9�����u������PS�5p���Y��YY������gu;�u������PS�5 p����Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�q�����0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u��y�������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF��0  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t����������������� Y���������������t������������������������� t
�������`p��������M�_^3�[葼���Ðyqzo�opTp_p�p�q��S��QQ�����U�k�l$���   �Pg3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|�����������uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�;�����h��  ��x���������>YYt�=px uV�r���Y��u�6����Y�M�_3�^�6�����]��[Ë�U��UV�uW��H�F��w�� �
�y�B��w�� ��t;�t�_+�^]Ë�U���S�u�M��b���3�9]u.�$��SSSSS�    �K�����8]�t�E��`p������   W�};�u+����SSSSS�    ������8]�t�E��`p������U�E�9XuW�u�:���YY�4V�E� �M�QP�����E����M�QP������G;�t;�t�+���^8]�t�M��ap�_[�Ë�U��V3�95lu09uu�U��VVVVV�    �|����������9ut�^]����V�u�u�������^]Ë�U���S3�VW9]��   �u�M��.���9]u.����SSSSS�    ������8]�t�E��`p������   �};�t˾���9uv(���SSSSS�    �������8]�t�E��`p����`�E�9Xu�uW�u��,  ��8]�tD�M��ap��;�E� �M�QP�^����E����M�QP�L�����G�Mt;�t;�t�+����3�_^[�Ë�U��V3�95lu99uu���VVVVV�    �8����������'9ut܁}���w�^]�H,  V�u�u�u������^]Ë�U��QSV��3�;�u���j^SSSSS�0����������   W9]w���j^SSSSS�0���������   3�9]���A9Mw	�f��j"�ЋM�����"w��]���9]t�-�N�E�   �؋�3��u��	v��W���0�A�E�3�;�v�U9U�rڋE�;Er�럈I���I�G;�r�3�_^[�� ��U��}
�Eu
��}jj
�j �u�u�M�����]Ë�U���4S3��E�VW���]��]��E�   �]�t	�]��E��
�E�   �]��E�P�-  Y��tSSSSS�������M� �  ��u�� @ u9E�t�M������+ú   ��   �tGHt.Ht&�K������.��j^SSSSS�0�V������  �U����t��   u��E�   @��}��EjY+�t7+�t*+�t+�t��@u�9}����E���E�   ��E�   ��E�   ��]��E�   #¹   ;��   ;t0;�t,;�t=   ��   =   �@����E�   �/�E�   �&�E�   �=   t=   t`;������E�   �E�E�   ��t�p���#M��x�E�   �@t�M�   �M�   �M��   t	}�� t�M�   ��E�   릨t�M�   �Y�������u������������    �   �E�=@�S�u��    �u�E�P�u��u��u�׉E���um�M��   �#�;�u+�Et%�e����S�u�E��u�P�u��u��u�׉E���u4�6������@������D0� ��L�P�S��Y�'��� �u  �u����;�uD�6������@������D0� ��L���V���Y�u�� �;�u������    룃�u�M�@�	��u�M��u��6�������Ѓ�����@�Y��Y�M����L��Ѓ�����@����D$� ��M��e�H�M���   �����  �Etrj���W�6�J�����E�;�u�N���8�   tN�6�ON�������j�E�P�6�]���������uf�}�u�E�RP�6��'  ��;�t�SS�6�6J����;�t��E���0  � @ � @  �}u�E�#�u	M�	E�E#�;�tD=   t)= @ t"=   t)= @ t"=   t= @ u�E���M�  #�;�u	�E���]��E   ��  �E�@�]���  �E��   �#�=   @��   =   �tw;���  �E�;��y  ��v��v0���f  �E�3�H�&  H�R  �E���  �E�   �  jSS�6� ������t�SSS�6����#���������j�E�P�6�5���������t�����tk����   �}�﻿ uY�E���   �E�;���   ���b������P���jSS�6��������C���SSS�6������#����   �����E�%��  =��  u�6�DL��Y���j^�0���d  =��  uSj�6�HH�������������E��ASS�6�-H������E�﻿ �E�   �E�+�P�D=�P�6�B������������9}�ۋ������@������D$�2M���0�������@������D$�M�������
ʈ8]�u!�Et��ȃ�����@����D� �}��   ���#�;�u|�Etv�u�� �S�u�E�jP�u������W�u�@����u4�L�P�����ȃ�����@����D� ��6����Y�����6������@��������_^[��jh�Q��0��3��u�3��};���;�u���j_�8VVVVV誼�������Y��3�9u��;�t�9ut�E%������@tu��u�u�u�u�E�P���i������E��E������   �E�;�t���0���3��}9u�t(9u�t�����������@��D� ��7�3���YË�U��j�u�u�u�u�u������]Ë�U���SV3�3�W9u��   �];�u"���VVVVV�    轻���������   �};�t��u�M�虯���E�9pu?�f��Ar	f��Zw�� ���f��Ar	f��Zw�� CCGG�M��tBf��t=f;�t��6�E�P�P�%  ���E�P�P�u%  ��CCGG�M��t
f��tf;�t�����+��}� t�M��ap�_^[�Ë�U��V3�W95lu3�9u��   �};�u���VVVVV�    �Ϻ���������`�U;�t��f��Ar	f��Zw�� ���f��Ar	f��Zw�� GGBB�M��t
f;�tf;�t�����+��V�u�u�u�w�����_^]Ë�U��} u3�]ËU�M�Mt�f��tf;uAABB����
+�]Ë�U����  ��f9Eu�e� �e�   f9Es�E��gf�Af#E���E��@�u�M��ܭ���E��p�p�E�Pj�EP�E�jP�$  ����u!E��}� t�E�`p��E��M#��Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5hzN�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�dz��+hz;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5hzN�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��lzA����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;`z�lz��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�`z�tz�3�@�   �tz�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+lz��M���Ɂ�   �ًpz]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�zN�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�|z��+�z;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�zN�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���zA����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;xz��z��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�xz��z�3�@�   ��z�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+�z��M���Ɂ�   �ً�z]���@u�M�U�Y��
�� u�M�_[�Ë�U���|�Pg3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u���SSSSS�    踮����3��O  �U�U��< t<	t<
t<uB��0�B���/  �$�1��Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �#  =�����/  � {��`�E�;���  }�ع`|�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9U�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �;����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[�͛�����W�����%�]�q�̕��6�+�ڕ��U���t�Pg3ŉE�S�]VW�u�}�f��E��U�� �  #��E��A�#�f�}� �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   t�C-��C �u�}�f��u1��u-��u)3�f9M�f�����$ �C�C�C0�C 3�@�  f;���   3�@f��   �;�u��t��   @uh��Sf�}� t��   �u��u;h��;�u0��u,h��CjP趝����3���tVVVVV�ʥ�����C�*h��CjP芝����3���tVVVVV螥�����C3��s  �ʋ�i�M  �������Ck�M��������3���f�M� {�ۃ�`�E�f�U�u�}�M�����  }�`|�ۃ�`�E�����  �E�T�˃������h  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��z����M�����?  ��  f;���  �]��E�3��ɉU��U��U�U��U�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��U���3�3�f9u���H%   � ���E��[���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �_�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[賒���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95����  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E������Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��3�PPjPjh   @h��D���zá�zV�5 ����t���tP�֡�z���t���tP��^áPg��3�9������Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v�����j^SSSSS�0�	��������V�u�M������E�9X��   f�E��   f;�v6;�t;�vWSV����������� *   ����� 8]�t�M��ap�_^[��;�t2;�w,�c���j"^SSSSS�0苙����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�h�;�t9]�^����M;�t����L���z�D���;��g���;��_���WSV�������O�����U��j �u�u�u�u�|�����]�U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U���SVW3�jSS�u�]��]��[����E�#��U���tYjSS�u�?�����#ʃ����tA�u�}+����   ;���   �   Sj�L�P�`��E���u�����    ����� _^[��h �  �u�  YY�E���|
;�r�����P�u��u�
�������t6�+��xӅ�wϋu��u��u��   YY�u�j �L�P�P�3��   �G����8u�*����    ����u��;�q|;�skS�u�u�u�D���#�����D����u�-���YP�H������H��E�#U���u)������    ��������L���u�#u��������S�u��u��u�٫��#���������3��������U��S�]V�u������@�������0�A$�W�y����   ���� @  tP�� �  tB��   t&��   t��   u=�I��
�L1$��⁀���'�I��
�L1$��₀���a��I��
�L1$�!���_^[u� �  ]����% �   @  ]Ë�U��EV3�;�u����VVVVV�    �ڕ����jX�
���3�^]Ë�U����  �ȃ�f9M��   S�u�M�蛉���M�Q3�;�u�E�H�f��w�� ���aV�   ��f9u^s)�E�Pj�u�9��������Et9�M싉�   f����q�M�jQj�MQPR�E�P�*  �� ���Et�E�8]�t�M�ap�[�Ë�U����u�M�������}�}3���u�u�u�u���}� t�M��ap��Ë�U����Pg3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[聆���Ë�U����u�M������E��~�M��Jf�9 t	AA��u���+�H�u �uP�u�u�u�p��}� t�M��ap����%0������̋M�������M����m����T$�B�J�3��������%镂���M������M����?����T$�B�J�3��ʅ����%�g����M���(���M��$`���M��`���M���(���M���(���M��`���M���_���M���_��h�h�   h ~�E�P�L����ËT$�B�J�3��S���� &������M��(����l����z(���M��r(���M���s���M��_���M��Z(���M��_���M��J(����l����?(����4����4(����P����)(���M��!(���M��I_���M��A_���M��9_���M��1_���M��)_���M���'���M��_���M��_���M��	_���M��_���M���^���M���^���T$�B��0���3��i�����&�����M���r���M���^���M��'���T$�B�J�3��6�����'�Ӏ���M��^��h�h�   h ~�EP��J�����h�h�   h ~��H���P�J����ÍM��U^���M��M^���E����   �e���M��5^��ÍM��,^���M��$^���T$�B��D���3�蜃����'�9��������̍M���]���E����   �e���M��]��ËT$�B�J�3��Z����H(�������̍M��v���M��Ј���T$�B�J�3��+����|(�����M���u���M�饈���E����   �e���M�m]��ËT$�B�J�3�������(����M��u���M��a����T$�B�J�3�輂����(�Y���M��nu���E����   �e���M��&���ËT$�B�J�3�耂��� )����M��2u���M�������T$�B�J�3��U����T)��~���M��u���M��χ���E����   �e���M�g%��ËT$�B�J�3�������)�~���M�s\���T$�B�J�3�������)�~���M��P\���T$�B�J�3��ˁ����)�h~���E����   �e���M�\��ÍM��\���M��\���M��\����p�����[���M���[����P�����[���M���[���M���[���M���[����`�����[����@����[���M��[���T$�B��@���3��(����*��}���M������M��������M���0�����M���H�����M���`�~����M���x�s����M����   �e����M����   �W����T$�B�J�3�貀����*�O}���M��4����M����)����M���0�����M���H�����M���`�����M���x������M����   ������M����   ������T$�B�J�3��<�����*��|���M��Z����|����Z��������Z����<����}Z���M��uZ���M��mZ���M��eZ����\����ZZ���M��RZ���M��JZ����L����?Z����l����4Z����,����)Z���������Z���������Z��������Z����������Y����������Y���M���Y���M���Y����l�����Y����L�����Y���M���Y���T$�B������3��<���`+��{���������Y��������Y���������Y����(����zY���M��rY���������gY����x����\Y���������QY���������FY����(����;Y��������0Y���������%Y����x����Y����H����Y����H����Y����h�����X����X�����X����x�����X����������X���M���X����������X����X����X����h����X���������X���������X���������X���������X��������xX���������mX���������bX���������WX����h����LX���M��DX���M��<X��������1X����x����&X���������X���������X���������X����������W���������W����8�����W����X�����W����h�����W���M���W���M��W����(����W����H����W����8����W���������W���������W���������|W���������qW���������fW��������[W����8����PW����X����EW���M��=W���M��5W���������*W���������W����8����W���T$�B��T���3��|���\,�)y���M���V����\��������0�������M���V���M���V���M���V����0�������M��V���M��V���M��V���M��V���M��V���M��V���M��}V���M��uV���M��mV���M��eV���M��]V���M��UV����L����JV����x����?V���M��7V���M��/V���� ����$V���� ����V��������V���M��V����<�����U���M���U����h�����U���M���U���M���U���M���U���� �����U����<����U����h����U���T$�B������3��'{����.��w���M�U����P����~U���M��vU���M��nU���M��fU����`����[U����|����PU���M��HU����@����=U���������2U��������'U��������U����$����U���������U����4��������M������M������p�������M���T���M���T���M���T����|����T���M��T���M��T����|����T���T$�B������3��z����/�v���M��L���M��tT���M��lT����D����1����D����&���M��NT���M��FT���M��>����M��6T����p����+T���M��#T����P����T����4����T���M��T����`�����S���M���S���M���S���T$�B��0���3��by����0��u������������M��S���M��S����t����v����t����k���� ����S����8����U���M��}S���M��uS����t����:����t����/���������$���M��LS���M��DS����t����	����t��������M��&S���M��S���M��S���M�������M������M���R���M���R���M���R���M���R���M���R���M���R���M���R���M���R���M��R���������R���������R���������R���M������� ����R���M��R���M��zR���M��rR���������gR���������\R���������QR���M��IR���M��AR���������6R���������+R��������� R���������R����t����
R����t�����x����������Q����\�����Q���M���Q���M���Q��������龳����������Q���M��Q����t����Q����\����Q���M��Q���M��Q����t����Q����\����Q���������tQ���T$�B��P���3���v���t1�s�������̋E����   �e���M�8Q��ËT$�B�J�3��v����3�Os�������������̋E����   �e���M����ËT$�B�J�3��rv����3�s�������������̍M��P���M�鰲���T$�B�J�3��;v����3��r���M�鍲���M��e���T$�B�J�3��v���,4�r���M��rP���M��h���M��{���M��h���M��r{���M��:����M�����T$�B�J�3��u���P4�Zr���M��P���M��gh���M��/{���M��Wh���M��{���M������M�����T$�B�J�3��ju����4�r���M���O���M��h���M���z���M��h���M���z���M�锱���M���g���M��z���M��\���T$�B�J�3��u���5�q���M��iO���M��g���M��yz���M��g���M��iz���M��1����M��	���T$�B�J�3��t���t5�Qq����0����O����0����O����������N����������N����������N����@�����N����������N����������N���������N�������� x���T$�B��p���3��(t���J�3��t����5�p���M��N���T$�B�J�3���s���L6�p���M������M���$�"���M���@����M���\����M����   �N����T$�B�J�3��s���p6�Fp���M��k����M��$�����M��@�����M��\����M���   ������M���   �q���T$�B�J�3��Is����6��o�������������������M����x����M����h����M����0����|M���� ����qM����@����fM����h����[M����x����PM����@����EM���� ����:M����0����/M����x����$M��������M���� ����M����d����s�����T�����L����h�����L����x�����L����@�����L���� �����L����0�����L����h����L����x����L����@����L���� ����L����0����L����x����L����h����tL����P����iL��������^L���� ����SL����P����HL���������=L���������2L���T$�B������3��q���J�3��q���7�=n���E���   �e���M�ҁ��ÍM��YN���M��QN���T$�B�J�3��\q���d8��m���������+����������K����p����K���������K���������K���������K���������yK����������M����P����M���������8�����������Q��������P�5��YÍ������4K��������P��4��YËT$�B������3��p���J�3��p����8�1m���������Ӏ���������Ȁ���������M�����������J���������J����t����J����@����J����(����J��������J����t����J���������J����(����zJ����@����oJ����l����dJ���������YJ����P��������P��������t����8J����P����L����l����rL����������P���������J����P����qL����l����FL���������P����8���� ����� ����������T��������T�������T$�B��L���3��7o���J�3��-o���$9��k���������I���������I���������vI���������kI���������0���������%���������JI���������?I����������������������������~���������I���������I����������H����������H����������H����d�����H����������H����������H����d����H���������H���������H���������H����t����H���������H����T����yH����D����nH���T$�B������3���m���J�3���m���@:�yj�������̋M��8H���M����   �*H���M����   �H���M����   �H���T$�B�J�3��m���\;�&j����̋M���G���M����   ��G���M����   ��G���M����   �G���T$�B�J�3��9m����;��i����̋M����d���T$�B�J�3��m��� <�i�����������̋M���H�(���T$�B�J�3���l���L<�}i�����������̋T$�B�J�3��l����<�Xi������̋EP�M�Q�]����ËT$�B�J�3��l���8=�'i�����̋M��H4���T$�B�J�3��cl���d=� i��������������̋EP�M�Q�S]����ËT$�B�J�3��*l����=��h�����̋M��_���M�����H���M��� ��H���M���<��H���M���X��H���T$�B�J�3���k����=�th��̋M��\_���M����H���M��� �H���M���<�H���M���X�|H���T$�B�J�3��k���4>�$h��̍M��XH���T$�B�J�3��ck���J�3��Yk����>��g����̍M��(H���T$�B�J�3��3k���J�3��)k����>��g����̋M��t���T$�B�J�3��k����>�g��������������̋EP��.��YËE����   �e���M��G��ËT$�B��\���3��j���?�Qg���������������̍M��xG���T$�B�J�3��j���J�3��yj���H?�g����̍M��HG���T$�B�J�3��Sj����?��f��������������̍M���]���T$�B�J�3��#j���@��f��������������̋E�P��-��YËE����   �e���M���F��ËT$�B��\���3���i���l@�qf���������������̋EP�M�Q��Z����ËT$�B�J�3��i����@�7f�����̍M��hF���M��`F����l����UF���T$�B��t���3��]i���A��e��������̋M��Mr���T$�B�J�3��3i����A��e��������������̋M���0���T$�B�J�3��i����A�e��������������̍M������T$�B�J�3���h����A�pe��������������̋T$�B��l���3��h���J�3��h���HB�;e���������̍�����%����P����%���T$�B��L���3��bh����B��d�������������̋EP�M�Q�SY����ËT$�B�J�3��*h���lC��d�����̋M���P�5#���T$�B�J�3�� h����C�d�����������̍M��$���T$�B�J�3���g����C�pd��������������̍M�X����T$�B�J�3��g����C�@d��������������̍M��hD���E�P�M�Q�X����ËT$�B�J�3��bg���J�3��Xg���XD��c���̍M������T$�B�J�3��3g����D��c��������������̋M��X9���T$�B�J�3��g����D�c��������������̋E����   �e���M��X��!��ËM����!���T$�B�J�3��f���8E�Qc���������������̋E����   �e���M��P�!��ËM���!���T$�B�J�3��df���tE�c���������������̍M��8���T$�B�J�3��3f����E��b��������������̍M��X8���M������T$�B�J�3���e���4F�b������̍M���B���M���B���T$�B�J�3���e���J�3���e����F�^b������������̋M����B���T$�B�J�3��e���4G�-b�����������̍M,�F���M�F���T$�B�J�3��[e���hG��a������̍M,�hF���M�`F���M��XF���T$�B�J�3��#e����G��a��������������̋M��(����T$�B�J�3���d����G�a���������������h�jh ~�E�P�{+����ÍM��/?���M��w����T$�B�J�3��d���H�?a�������������̋T$�B�J�3��{d���pH�a������̋M��:���T$�B�J�3��Sd����H��`��������������̋M��X����M���@齑���M���X鲑���T$�B�J�3��d��� I�`���E�P��'��YËT$�B�J�3���c���,I�`���M��mW���T$�B�J�3���c���XI�a`���M��F����T$�B�J�3��c����I�>`���M��#����M����h@���T$�B�J�3��sc����I�`���M���V���u��M'��YËT$�B�J�3��Fc����I��_���M��@���T$�B�J�3��#c���J��_���T$�B�J�3��c���M�_����hP�����Yù�~��U��h�������Y�h�������Yù@��U��h���چ��Y�h���Ά��YÃ=�} uK��}��t��}�Q<P�B�Ѓ���}    ��}��tV�����V�Z&������}    ^ù�~�U����~������@�U���A�]��                                                   dS rS �S �S �S �S T T $T @T XT pT �T �T �T �T �T �T 
U U ,U 8U FU \U nU zU �U �U �U �U �U �U �U V V  V *V :V DV PV bV vV �V �V �V �V �V �V �V �V  W W W .W BW NW `W vW �W �W �W �W �W X X *X DX PX bX tX �X �X �X �X �X �X Y  Y 0Y @Y RY `Y nY ~Y     �S         �.�D� �"�        �Y͙d�����        �3�                    ΁qP       ~   � �� bad allocation   �$ � �  � !  ��    @u3D-COAT     c:\program files\maxon\cinema 4d r12\plugins\applink_cinema4d\source\applinkdialog.cpp  Start import!   To import a new object? File exists!    export.txt  Folder ..\MyDocuments\3D-CoatV3\Exchange not found! 3D-CoatV3   Exchange    preference.ini  3D-Coat.exe is run! 3D-Coat.exe not found!  open                c:\program files\maxon\cinema 4d r12\plugins\applink_cinema4d\source\applinkexporter.cpp    
   c:\program files\maxon\cinema 4d r12\resource\_api\ge_dynamicarray.h    ]   autopo  curv    prim    alpha   vox retopo  ref uv  ptex    mv  ppp [   # end   v       # begin      vertices
            �?vt   texture vertices
  /   f   usemtl   faces
 g   mtllib  mtl map_    illum 2
    Tr 0.000000
    Ns 50.000000
   Ks  Kd  Ka 0.300000 0.300000 0.300000
  newmtl  No selected objects!    Object "    " has no UVW tag.
UV coordinates can't be exported. Material not found on   object. Default Name    Export object   #Cinema4D Version:  %d.%m.%Y  %H:%M:%S  #File created:  #Wavefront OBJ Export for 3D-Coat
  File     write success! [SkipExport]
   [SkipImport]
         �import.txt  output.obj  obj �p� ? ���� T�8�� L��  � �� P� 0� �� �� �� �  � @�       Y@�0 �  � �  � �� 0� �p	�� �� P� � `� ���
 � � P� �� 0� �p	�� P� � `� 0��  �  � 00PpSelection   Error on inserting phongTag. Object:    Create objects...   Memory allocation error for material.   ���4 &��  @0� �p	�)�*P`�@$0#�pP%��0#�P%�vector<T> too long  bad cast    ios_base::eofbit set    ios_base::failbit set   ios_base::badbit set    \ G    X       P    can not removed!   normalmap   displacement %f displacement    map_Ks %s   map_Ks  map_Kd %s   map_Kd  Ke %lf %lf %lf  Ke  Ks %lf %lf %lf  Ks  Ka %lf %lf %lf  Ka  Kd %lf %lf %lf  Kd  illum %d    illum   d %lf   d   Ns %lf  Ns  newmtl %s   Open file   .    not found!     c:\program files\maxon\cinema 4d r12\plugins\applink_cinema4d\source\applinkimporter.cpp    Wrong face in OBJ file! f   vt  Gathering of data...        �dy���=vt %lf %lf %lf  vt %lf %lf  v %lf %lf %lf   g %s    mtllib %s   Parse file...   Open file:  textures.txt     �[�Y��@���P�p�`�icon_coat.tif   c:\program files\maxon\cinema 4d r12\plugins\applink_cinema4d\source\applinkpreferences.cpp pPPPPPP0\          �?��c�n�o`i0e�e0j     �f@-DT�!	@ �Р� �� �0��@u     @�@ �Р� �� �0��0�d������@�P����`�0�p�P�c:\program files\maxon\cinema 4d r12\resource\_api\c4d_gui.cpp  � �Р� �� �0��`�� �Р� �� �0�� �����������о���0�@�� �Progress Thread 0%  ~   %       c:\program files\maxon\cinema 4d r12\resource\_api\c4d_file.cpp c:\program files\maxon\cinema 4d r12\resource\_api\c4d_general.h    %s         ����MbP?| �� p� `�    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_baseobject.cpp   c:\program files\maxon\cinema 4d r12\resource\_api\c4d_resource.cpp #   M_EDITOR    ! �res c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basetime.cpp      �Ngm��C   ����A  4&�k�  4&�kC$!�� PP    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_pmain.cpp        �������������c:\program files\maxon\cinema 4d r12\resource\_api\c4d_libs\lib_ngon.cpp        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basebitmap.cpp   l!�c:\program files\maxon\cinema 4d r12\resource\_api\c4d_gv\ge_mtools.cpp �!��!`H"�"�+*   C   �����";/�string too long invalid string position r            
   !   "   2   *            #   3   +       w   a   r b     w b     a b     r +     w +     a +     r + b   w + b   a + b   ,#6z:����t#n??Unknown exception   �#�??csm�               �                              �?      �?3      3            �      0C       �       ��                                                                                                                                                                                                                                                                                                        ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������LC_TIME LC_NUMERIC  LC_MONETARY LC_CTYPE    LC_COLLATE  LC_ALL  H�    !<�xm!0�xm�a$�xmY�xm�xmC	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ _., _   ;   =   =;  l�#w}?bad exception   EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    ��e+000          �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:    CorExitProcess  m s c o r e e . d l l         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow         �������             ��      �@      �              �?5�h!���>@�������             ��      �@      �        HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun united-states   united-kingdom  trinidad & tobago   south-korea south-africa    south korea south africa    slovak  puerto-rico pr-china    pr china    nz  new-zealand hong-kong   holland great britain   england czech   china   britain america usa us  uk  swiss   swedish-finland spanish-venezuela   spanish-uruguay spanish-puerto rico spanish-peru    spanish-paraguay    spanish-panama  spanish-nicaragua   spanish-modern  spanish-mexican spanish-honduras    spanish-guatemala   spanish-el salvador spanish-ecuador spanish-dominican republic  spanish-costa rica  spanish-colombia    spanish-chile   spanish-bolivia spanish-argentina   portuguese-brazilian    norwegian-nynorsk   norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg   german-lichtenstein german-austrian french-swiss    french-luxembourg   french-canadian french-belgian  english-usa english-us  english-uk  english-trinidad y tobago   english-south africa    english-nz  english-jamaica english-ire english-caribbean   english-can english-belize  english-aus english-american    dutch-belgian   chinese-traditional chinese-singapore   chinese-simplified  chinese-hongkong    chinese chi chh canadian    belgian australian  american-english    american english    american    �	ENU �	ENU �	ENU �	ENA �	NLB �	ENC �	ZHH |	ZHI t	CHS `	ZHH L	CHS 8	ZHI $	CHT 	NLB  	ENU �ENA �ENL �ENC �ENB �ENI �ENJ �ENZ �ENS hENT \ENG PENU DENU 4FRB $FRC FRL  FRS �DEA �DEC �DEL �DES �ENI �ITS �NOR xNOR dNON LPTB 8ESS (ESB ESL ESO �ESC �ESD �ESF �ESE �ESG �ESH xESM hESN TESI DESA 0ESZ  ESR ESU �ESY �ESV �SVF �DES �ENG �ENU �ENU �USA �GBR �CHN �CZE �GBR �GBR �NLD xHKG lNZL hNZL \CHN PCHN DPRI <SVK ,ZAF  KOR ZAF KOR �TTO �GBR �GBR �USA �USA 6-0   OCP ACP Norwegian-Nynorsk   c c s   U T F - 8   U T F - 1 6 L E     U N I C O D E    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   ->* &   +   -   --  ++  ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        �xl`TH<4(��pT@ $� �����p���������0�������,��������������|pd\P8,����xT8�������`XL<  ���\@������GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    1#QNAN  1#INF   1#IND   1#SNAN  CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           Pg $b   RSDS�2����C����]1E~   C:\Program Files\MAXON\CINEMA 4D R12\plugins\Applink_Cinema4D\obj\Applink_3DCoatR12_Win32_Release.pdb               `           $0L    `       ����    @    `        ����    @   h           xL                @`�           ���    @`       ����    @   �\`        ����    @   �           ��                x`           $,    x`        ����    @              Xd,    �`       ����    @   H           ��,    �`       ����    @   �            �`�           ��    �`       ����    @   ��`       ����    @               08    �`        ����    @               ah           x��     a       ����    @   hLa              P   �           ���    La       ����    @   ��`              @   ��`              @                La�            �a`           p��,    �a       ����    @   `            �a�           ��    �a        ����    @   �            �a�           �    �a       ����    @   �            0bD           Tdd,    0b       ����    @   D    P       Pb�           ����     Pb       ����    @   �            �b�           ��    �b       ����    @   �            �b8           HT�    �b       ����    @   8             c�           ���     c       ����    @   �             c�           ��T�     c       ����    @   �            @c            0@��    @c       ����    @        X       �cp           ����     �c       ����    @   p           ���    �c       ����    @   ��c        ����    @              �                �c4           DT��    �c       ����    @   4             d�           ��     d        ����    @   �            <d�           ���    <d       ����    @   �             `h            td,           <HL    td       ����    @   ,            �dx           ��    �d        ����    @   x            �d�           ��L    �d       ����    @   �            �d             , �L    �d       ����    @               X `     e        ����    @   H             ,e�            � �     ,e        ����    @   �             De�            � � `     De       ����    @   �             �c            �e8!           H!P!    �e        ����    @   8!            �e�!           �!�!    �e        ����    @   �!            �e�!           �!�!    �e        ����    @   �!            �e"            ","`     �e       ����    @   "             f\"           l"t"     f        ����    @   \"            Lf�"           �"�",    Lf       ����    @   �"            |f�"            ##T�    |f       ����    @   �"            \g@#           P#X#    \g        ����    @   @#            \`�            dc�#           �#�#�    dc       ����    @   �#            h�#           �#$�    h       ����    @   �#�2 �3 � �E �F � !� �� � �� L� �� �� � /� k� �� ڳ ��  � �� 9� �� �� \� �� λ �� �� 9� y� �� ۿ .� �� �� 7� �� �� B� �� >� �� J� �� � b� �� �� � 0� a� �� �� � d� �� �� �� 4� h� �� �� � Q� �� �� �� � @� �� �� �� � H� �� �� �� 7� �� �� ��  � [� �� �� �� I� p� �� �� � '� J� x� �� �� ��                 �����    �"�   �%                       �����    �"�   �%                       "�	   D&                       ����<�    D�   L�   T�    \�    d�    l�    t�    |�"�   �&                       ������    ��   ư����ΰ   ְ   ް   �   �   ��   �	   �
   �	   �   �   �   �   �   '�   /�   7�   ?�   G�   O�   W�   _�   g�   o�   w�������    ��   ��"�   �'                       "�	   �'                       �����������   ������   #�   <�   D�����б����ر����x�    p�"�   8(                       ������    ��"�   l(                       �����    ۲   �"�   �(                       �����    '�"�   �(                       ����J�    R�"�   )                       ������    ��"�   D)                       ������    ��   ��"�   x)                       ������"�   �)                       �����"�   �)                       "�   0*                       ����;�    T�    \�    d�    l�    w�    �    ��    ��    ��    ��    ��    ��"�   �*                       ����޴    �   �   ��   �   �   �   +�"�    +                       ����T�    \�   g�   r�   }�   ��   ��   ��"�   �+                       ����ʵ    ҵ   ݵ   �   �   �   �    ������   ��	   �
   �   �   �   &�   1�   <�   G�   R�   ]�   h�   s�   ~�   ��   ��   ��   ��"�B   �,                       ����ʶ    ն   �   �   ��   ��   ��    ��������   ��	   	�
   �   �   *�   5�   @�   K�   V�   a�   l�   w�   ��   ��   ��   ��   ��   ��   ��   ̷   ׷   �   �   ��    �!   �   �#   $�$   ,�%   4�&   ?�'   J�(   U�)   `�*   k�+   v�,   ��-   ��.   ��   ��0   ��1   ��2   ��3   ȸ4   Ӹ5   ޸6   �7   ��8   ��9   
�:   �;    �   +�=   3�>   ;�?   F�@   Q�"�$   �.                       ����z�    ��   ��   ��   ��   ��   ��   ��   ù   ˹    ӹ
   ۹   �   �    �   ��   �   �   �    �   &�   1�   9�   A�   L�   W�   b�   j�   u�   }�   ��   ��   ��    ��!   ��"   ��"�   �/                       ����ߺ    �   �    �   ��   �   
�   �    �   (�	   3�
   >�   I�   T�   _�   j�   u�   }�   ��   ��   ��   ��   ��   ��   ��   û"�   �0                       �����    ��   ��   �    �    �    "�    *�   2�   :�	   E�
   M�   X�   c�   k�   v�   ~�"�?   �1                       ������    ��   ��   ��    ʼ    ռ    �   �   �   ��   �   �   �   $�   ,�   7�   B�   J�   R�   Z�   b�   j�   r�   z�   ��   ��   ��   ��   ��   ��   ��   ��   Ƚ   ӽ!   ۽"   �"   �$   ��%   ��&   	�'   �"   �)   '�*   /�+   :�,   E�"   P�.   [�"   f�0   q�1   |�0   ��3   ��4   ��5   ��0   ��0   ��0   ��0   ˾:   Ӿ;   ۾<   �   ����� �"�   �3                       ����`�"�   �3                       ������    ��"�   �3                       ����˿    ӿ"�   4                       "�   t4                       ������������   �   �   �   �   &�"�   �4                       ����I�����Q�   Y�   a�   i�   q�   y�"�	   ,5                       ������������   ��   ��   ��   ��   ��   ��   ��"�   �5                       �����������   �   �   �   '�   /�"�
   �5                       ����R�����]�����h�����s�   ~�������   ��   ��   ��������������"�   D6                       "�   �6                       �����    �   �   )�   4�"�   �6                       ����]�    e�   p�   {�   ��   ��"�#   47                       ������    ��   ��   ��   ��   ��   ��   
�   �    �	   +�
   6�   A�   L�   W�   b�   m�   x�   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �   �   �    (�!   3�����f�    �    ��"�   L8                       "�   �8                       ������    ��   ��   ��   ��   ��    ��    ��   �    �	   �
   �
   1�    #�    <�"�   H9                       ����r�    }�   ��   ��   ��   ��   ��   ��   ��   ��	   ��
   ��   ��   �   �   �   "�   -�   8�   C�   C�   N�   Y�   d�   o�   o�   z�   ��   ��   ��   ��"�   d:                       ������    ��������   ��   �����������   &�   1�����<�����G�
   R�
   ]�   h�   s�   ~�   ��
   ��   ��   ��   ��   ��
   ��   ��   ��   ��   ������0�    8�   F�   T�"�   <;                       ������    ��   ��   ��"�   �;                           `�     �;   �;�;    @`    ����       ��     \`    ����       �>������"�   <                       ���� �"�   D<                       @           Z@           �����    ����                  "�   �<   �<                           �<              p<@                        �<����        P�����    "�    =   =               ������"�   \=                       @           ,             �=����        ������    "�   �=   �=               "�   >                       ������    ��   ��   ��   	�"�   X>                       ����0�    8�   C�   N�   Y�������"�   �>                       ������"�   �>                       ������"�   �>                       �����    ������"�   ?                       ����`�"�   @?                           p    �?������"�   |?                          �?�?�;     c    ����    (   �-    �b    ����    (    -    c?    ,@������"�    @                          8@�;    dc    ����       F?������    ��������"�   T@                       @           I1             �@����        @�����    "�   �@   �@                   %    <A����p�����x�������"�    A                          LAhA�;    @c    ����    (   3     c    ����    (   �2������"�   �A                       ������"�   �A                       �����"�   �A                       @           v7@           g7����    ����    ����    ����    "�   (B   lB                             B            B@           D;@           B:"�    C   �B                             �B            �B����    ����    ����p�              ����{�@           �?             0C����        ������    "�   TC   @C               ������"�   �C                       �����"�   �C                       ����@�"�   �C                       @           �E            D����p�           x�        "�   8D   $D               @           �H            |D"�   �D   �D               ����������    ����                         ������"�   �D                       �����            ,�"�    E                       ����`�            |�"�   \E                       @           >N            �E"�   �E   �E               ������                                     @           	P            F"�   XF    F               ������    ��                                     @           �T@           �S"�   �F   �F                             �F            �F����    ����    �����              ���������P�"�   ,G                       ������    ��"�   XG                       ������    ��   ��"�   �G                       ������"�   �G                       ���� �����9�   A�"�   �G                       @           �k@           �k����    ����    ����    ����    "�   PH   �H                             @H            0H������"�   �H                       ������    ��   ��"�   �H                       ������"�   $I                       �����"�   PI                       ����B�"�   |I                       ����e�    m�"�   �I                       ������    ��"�   �I                       ������"�   J                           0/    LJ   \J�?�;    |f    ����    (   �/����    ����    ����    YC    ����    ����    ����    �D    ����    ����    ����    �E    ����    ����    ����    �F    ����    ����    ����    �H        QH����    ����    ����    �H    ����    ����    ����    �I    ����    ����    ����    �K    ����    ����    ����    ?M    ����    ����    ����    vN    ����    ����    ����ERVR    ����    ����    ����    �T    ����    ����    ����    Z    ����    ����    ����    ol    ����    ����    ����    �x        �x        �x    ����    ����    ����    �y    ����    ����    ����        �~�~����    ����    ������@           ������    ����                  �L"�   �L   �L                   ����    ����    ����    ΁    >�G�����    ����    ��������    ����    ����    ����N�R�    l}    �M   �M�;    h    ����       �    ����    ����    ����    =�����    L�����    ����    ����    ������    �����    ����    ����2�6�    ����    ����    ��������    ����    ����    ����    i�    ����    ����    ����    ƕ    ����    ����    ����    ��    ����    ����    ����ϛ�    ����    ����    ����    ��    ����    ����    ��������    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    c�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ;�    ����    ����    ����    �    ����    ����    ����    )    ����    ����    ����    Q    ����    ����    ����    �D    ����    ����    �����N�N    ����    ����    �����OP    ����    ����    ����    �P    ����    ����    ����    �W    ����    ����    ����    Y    ����    ����    ����    �]    ����    ����    ����    Y_        �^����    ����    ����m'm    ����    ����    ����    =�R         �S  � \S         �S T�                     dS rS �S �S �S �S T T $T @T XT pT �T �T �T �T �T �T 
U U ,U 8U FU \U nU zU �U �U �U �U �U �U �U V V  V *V :V DV PV bV vV �V �V �V �V �V �V �V �V  W W W .W BW NW `W vW �W �W �W �W �W X X *X DX PX bX tX �X �X �X �X �X �X Y  Y 0Y @Y RY `Y nY ~Y     �S     C CloseHandle EProcess32Next Module32First CProcess32First  � CreateToolhelp32Snapshot  KERNEL32.dll  ShellExecuteExA SHELL32.dll �InterlockedIncrement  �InterlockedDecrement  !Sleep �InitializeCriticalSection � DeleteCriticalSection � EnterCriticalSection  �LeaveCriticalSection  �RtlUnwind -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent ZRaiseException  �GetLastError  �HeapFree  � DeleteFileA �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �LCMapStringA  zWideCharToMultiByte MultiByteToWideChar �LCMapStringW  [GetCPInfo �GetModuleHandleW   GetProcAddress  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �SetLastError  RGetACP  GetOEMCP  �IsValidCodePage �GetModuleHandleA  �HeapCreate  �HeapDestroy WVirtualFree TVirtualAlloc  �HeapReAlloc �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA �WriteFile �GetConsoleCP  �GetConsoleMode  AFlushFileBuffers  hReadFile  �SetFilePointer  �GetModuleFileNameA  ExitProcess JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW �GetEnvironmentStringsW  TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �HeapSize  �GetLocaleInfoA  =GetStringTypeA  @GetStringTypeW  mGetUserDefaultLCID  � EnumSystemLocalesA  �IsValidLocale �InitializeCriticalSectionAndSpinCount �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW �SetStdHandle  �LoadLibraryA  �GetLocaleInfoW   CreateFileW x CreateFileA �SetEndOfFile  #GetProcessHeap      ΁qP    �Y          �Y �Y �Y �� �Y   Applink_3DCoatR12.cdl c4d_main                                ��D�    .?AVApplinkDialog@@ D�    .?AVGeDialog@@  ����D�    .?AVbad_alloc@std@@ D�    .?AVexception@std@@ D�    .?AVfacet@locale@std@@  D�    .?AVcodecvt_base@std@@  D�    .?AUctype_base@std@@    D�    .?AVios_base@std@@  D�    .?AV?$_Iosb@H@std@@ D�    .?AV?$basic_istream@DU?$char_traits@D@std@@@std@@   D�    .?AV?$basic_ios@DU?$char_traits@D@std@@@std@@   D�    .?AV?$ctype@D@std@@ D�    .?AV?$basic_streambuf@DU?$char_traits@D@std@@@std@@     D�    .?AV?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    D�    .?AV?$codecvt@DDH@std@@ D�    .?AV?$basic_istringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    D�    .?AV?$basic_filebuf@DU?$char_traits@D@std@@@std@@   D�    .?AVlogic_error@std@@   D�    .?AVruntime_error@std@@ D�    .?AVlength_error@std@@  D�    .?AVfailure@ios_base@std@@  D�    .?AVbad_cast@std@@  D�    .?AV?$basic_ifstream@DU?$char_traits@D@std@@@std@@  ����D�    .?AVCommandData@@   D�    .?AVBaseData@@  D�    .?AVApplinkPreferences@@    ��D�    .?AVTriangulator@@  D�    .?AVCTriangulator@TRIANGULATOR@@    ������D�    .?AVGeModalDialog@@ D�    .?AVGeUserArea@@    D�    .?AVSubDialog@@ D�    .?AViCustomGui@@    ����������������������D�    .?AVGeSortAndSearch@@   D�    .?AVNeighbor@@  D�    .?AVDisjointNgonMesh@@  ����������������D�    .?AVC4DThread@@ ������������������D�    .?AVGeToolNode2D@@  D�    .?AVGeToolDynArray@@    D�    .?AVGeToolDynArraySort@@    D�    .?AVGeToolList2D@@  ����������D�    .?AV_Locimp@locale@std@@    ��   ��D�    .?AVout_of_range@std@@  ������������ � ���� �(�0�8�        ��
   Copyright (c) 1992-2004 by P.J. Plauger, licensed by Dinkumware, Ltd. ALL RIGHTS RESERVED.              N�@���D��D�    .?AVtype_info@@             u�  s�          ��            fmod         TZv��v���v��v���7��v�v��v�sqrt    �
�   �        ��D�    .?AVbad_exception@std@@ ��������    ��                                                                                                                                                                                                                                                                                                                                                abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     Ph�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����    C                                                                                              xm            xm            xm            xm            xm                              w        ����Pv�m   �mPh                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                         �M�M�M�M�M�M�M�M�M�M                                                                                                                                                                                                                                                                                         `�    `�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����
                                                             0   	   � 
   @        ��   ��   ��   \�   4�   ��   ��   ��   |�   �    ��!   ��"   H�x   4�y   $�z   ��   ��    ���      x   
   ?         ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      �����������������������)�.�J�Z�n�~��������������"�B�G�a�f��������������
�*�>�V�j��������������� . 3 M R r � � � � � � � *B  ������������|plhd`\XTPLHD@8,$\���������	         Pv.   w؈؈؈؈؈؈؈؈؈w   .       �                                                                                                                                                                                                                                   �&             $         �   �!   �         �   �   �   �   �    �   �   �   �   �   �   �   �   �   �"   �#   �$   �%   �&   �      �      ���������              �       �D        � 0     �    �p     ����    PST                                                             PDT                                                             �y z����        ����           ���5      @   �  �   ����             ������������   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l           �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                       �   0040E0q0�0�0�0�0�0�0f1t1�1�1�1�1J243]3�3�3�3P4f4}4�4�4�4�45%565N5v5�5�5�5�7�7�7�899-9E9R9�9:,:A:Z:g:�:�:�:�:�:�:�:;!;5;I;\;j;�;�;<j<�<�<�< =6=L=�=�=�=>F>s>�>�>?=?�?�?�?      �   &070�011]1o1�1�1�1�1<2F2�2�2�2�2�2(3S3e3u3�3�3�3�3414K4d4$7V7g7�7�7�7�78858\8u8�8�8�8�8U9s9�9�9�9:(:�:�:�:�:�:�:;;F;W;�;�;�;6<G<�<�<�<=F=W=�=�=>V>g>�>�>?V?f?w?�?�?�?�?   0  �   &080I0[0n0z0�0�0�0�0�1�1�1�1�1�1�1252]2}2�2�2�23(3E3e33�3�3�344I4^4p4�4�4�4�4�4�4�4�4�4�4 55555&565f7v7�8�8�899999N9�9�9�9�9�9:I:[:m:v:�:�:�:�:�:�:�:;<&<?<X<p<�<�<�<�<�<==3=H=a=|=�=�=�=�=�=>M>c>y>�>�>�>�>�>?V?k?�?�?�?�?�?�?   @    30L0e0}0�0�0�0�011)1>1G1`1u1}1�1�1�2�2 3313J3c3~3�3�3�3�3�34.4K4l4�4�4�4�4�4�4�4�45555T6j6�6�6�6�6�67737K7d7}7�7�7�7�7�788.8@8I8_8q8y8�8�8�9�9�9:):B:[:v:�:�:�:�:�:; ;;;i;z;�;�;�;�;�;�;�;�;<,<J=`=y=�=�=�=�=�=>)>A>Z>s>�>�>�>�>???5?G?�?�?�?�?�?   P  ,  0 0;0_0�0�0�0�0�01�1�1�1�1�1�122!232�2�2�2�2�23,3;3s3�3�3�3�3�3�34!474M4b4x4�4�4�455!535t5�5�5�5�5�5�5646O6d6m6�6�6�6�6777I7[7d7y7�7�7�7�78(8:8X8w8�8�8�8�8�8!939E9Q9f99�9�9�9:':9:D:Y:r:�:�:�:;!;3;?;T;m;�;�;�;�;�;<<-<w<�<�<�<�<�<==B=[=t=�=�=�=�=>0>_>p>�>�>�>�>�>�>�>�?�?�?   `  �   0-0F0_0w0�0�0�0�0�01!1�1�1�1�12 2V2l2�2�2�2�2�2�2333J3c3x3�3�3�3�364K4f4�4�4&585J5f5�5/6C6\6q6z6�6�6�6�67757J7f7�7�7�7�7�7�7�78D8[8j8�8�8�8�8�89999U9p9�9�9�9�9�9�9:":4:F:N:h:�:�:�:F;[;�;<<c<x<�<�<�<7=M=e=�=>>6>�>�>�>?h?�?�?   p  �   Y0�0�0�01(1A1Q1�1�1�1�1�1%272c2�2�2�23373M3�3�3�34}4�4�4�45'5@5V5�5�5�56646L6b6�6�6�67&7;7O7Z7�7�7�7�7�7	8=8V8{8�8E9�9�9�96:j:�:�:�:�:�:;;I;�;�;�;D<`<|<�<h=   �  p   j1�1�25I5�5�5�5�576O6h6}6�6�677"787I7T7�7�7�7�7	8?8e8z8�8�8�8A9":0:�:;�;�;"<0<�<�<i=y=�=�=@>N> ?
?&? �  �   �0�0�002>2�2�23B4L4o465D5\5t5�5�5b6x6�7V8e8�8�8969H9�9�9�9�9�9":D:g:�:�:�:D;�;�;6<H<^<p<�<�<�<=�=�=>A>l>�>�>??0?B?�?�?�?   �  �   @0�0�0
1K1�1�1�1�1�1282b2�2)3^3�3�34D4�4�4�4�4�4585b5�5)6o6�6�67(7a7�7�7�78�8�89�9�9�9�9�9:b<�<�<�<==G=`=�=�=�=>8>�>�>)?Q?f?�?�?�?�?�? �  �   b0�0�0�0[1�1�2�2o3�3/4@4R4k4�4�4Q5�5�5�5�6�6717A7P7�7�7�7�78"8z8�8�8�8�8�8.9C9X9m9u9�9�9�9:,:I:^:�:-;9;N;�;�;<Y<u<�<�<!===~=�=�=�=8>T>�>�>�>%?G?�?   �  �   00J0Z0i0�0�011&1;1�1�1�1�1�12>2P2�2�2�2�2�2?3W3p3�3�304E4�4�4 5u5�5�5!6>6j6�6�6(7>7�7z8�8�8�8�8�8�8�8U9m9�9�9�9�9::�:�:�;�;X<m<�<�<�<�<�<�<5=N=g==�=�=�=�=>'>�>�>W?   �  �   �0�2�2�2�2�23�3>5v5�5$696M6U6n6�6�6�6�6707H7a7�7�7�7�7�788(8A8�8�8�8�8�89;9Z9m9�9:5:�:�:c<w<�<�<"=�=5>?>p>�>�>�>?A?c?�?   �  �   c12�4�5&6�6B7x7f8x8�8�8�8�8989O9h9�9�9:$:\:�:�:�:U;v;�;�;<<-<A<�<�<�<�<�<0=N=b=k=�=�=�=> >8>Q>�>??!?:?N?W?o?�?�? �  t   0040�01*162D2Z2�2�2�2�23$3:3V3o3�3�3�3�5�5�5�5v6�6�6�6�6�6	7"7i8t8�8�8)949�9�9�9�9}:�:�:�:�;�=�=�=�>�>     <   %0�0�001�12
2<2�2�2>4I45525�6::2:D:R:|:�>�?�?    0   u02(2�2%3�3�3�3�4�4u5�5�5V6f6F:U:&>5>     \   '2�2�2�2!383�3�3�364K45X5&656Y:2;�<�<�<�<
==&=5=\=�=�=�=�=�=>>>>+>}>�>�>?*?�? 0 `   �0�0�1�1�1222;2F2P2v2�2�2�2�2!3�3�34%4<4^4�4�4�5�5�8�8�=�=>>7>?>E>J>[>�>�>�>v?�?   @ T   &040Q0p0�0�1�133}3�45�557f7x7�8F:T:;;9;@;V;�;�;�;<<9<@<V<�<�<�<j>�>�> P L   5062E2�5�5�7�7�8�8d9�9�9�9�9:':8:?:i:�:�:�:6;D;j;�;�;"<<<�=F?�?�?�? `    0F0S01�2�2f:x:6=D= p �   �1�1�1�1�12$2D2a2t2�2�2�23$3T3�3�3�3�34�4�4 55D5�5�5�6�6�6�6�6�67A7a7�7�78 8�8�8�89<9z9�9�9�9:[:�:�:$;`;�;�;<1<L<e<~<�<�<�<==j=�=�=�=�=�=6>c>u>�>�>�>?5?[?�?�?�?�?   � �   	060H0�051=1�1�1;2�2�23=3h3�3�34I4c4�4�45K5v5�5�56.6T6�67�7�7%8d8�8�8�8=9�9�9:a:�:�:�:2;k;�;�;�;�;�;1<j<�<�<t=�=>`>�>�>@?�?�? � |   S0�01S1�12s2�233�3�3S4�45c5�5#6�6�67�7�7@8p8�8�8 909`9�9�9 :M:q:�:�:�:;N;�;�;
<[<�<�<>=~=�=�=">D>�>�>�>$?d?�?�? � �   050N0t0�0E1J1U1k1�1�1242n2@3�344 4$4(4,4044484f45p5t5x5|5�5�5�5�5�566X6b6�6�6�6�67!7A7a7�7�7�78$8D8t8�8�8$9D9t9�9�9�9�:�:�:;$;T;�;�;�;	<&<8<J<h<�<�<�<�<�<�<=!=5=S=l=~=�=�=�=�=�=>d>�>�>�>?D?�?�? � �   0T0l0�0�01T1�1�1�1�2�2�23.3U3�34484R4'5d5�5�5�56686B6d6�67$7D7f7z7�7�7�7S8�8%9y9�9�9:4:a:�:C;s;�;�;�;<A<V<j<<�<�<=Q=�=�=�=�=�=�=$>T>Q?�?�?�?�?   � �   0050p0�0�0�0�0�0:1^1w1�1�12!222Y2�2�2�2�2�233?3_3}3�3�3�34P4�4�45�5�5�5$6S6}6�6�6�627d7�7�7�788-8I8W8w8�8�8�8�8�899/9D9_9q9�9�9�9�9�9�9�;�<�<=d=�=9>�>�>4?U?�?�? � �   t0�0H1i12-2V2i2{2�2�2�2�2363i3�3�3�344_4q4�4�4�4�45=5K5[5�6�677k7�7�7�78$8Q8b8�8�8�8�8�8�899#9A9R9t9�9�9�9�9::0:@:d:�:�:�:�:�:�:;;0;?;O;`;�;�;�;�;�;<4<T<t<�<�<�<�<�<$=D=t=�=�=�=�=>$>T>q>�>�>�>�>?!?1?A?T?t?�?�?�?�?   � (  040T0t0�0�0�0�011,1�1�1�1252t2�2�2�2�2343T3t3�3�3�3�34!444a4t4�4�4�4�4�4�45!505Q5t5�5�5�5�5�566$6D6_6m6{6�6�6�6�67$7D7d7�7�7�7�7808A8]8�8�8�8�8�8�8$9D9d9�9�9�9�9�9::.:@:d:~:�:�:�:�:�:;.;E;\;m;{;�;�;�;�;�;<&<5<E<V<�<�<�<�<==4=T=t=�=�=�=�=>4>T>t>�>�>�>�>?4?T?t?�?�?�?�?   � �   0D0p0�0�0�0�0141T1t1�1�1�1�1242T2t2�2�2�2�2343T3t3�3�3�3�34$4D4a4t4�4�4�4�4�45&5:5J5t5�5�5�5�5�5 656�6�6�6747T7q7�7�7Y8u8�8�8Y9u9�9�9:<:X:t:�:�:;5;�;<1<�<�<�<�<=4=A=o=�=�=�=�=>$>Q>d>�>�>�>�>?2?Q?t?�?�?�?   �   $0D0a0�0�0�0�01D1q1�1�1�12A2a2�2�2�2�23$3D3d3�3�3�3�3�3444T4�4�4�4l5�5�56q6�6
7-7�7�7�7a8~8�89.9C9�9�9:A:d:�:S;|;�;#<L<t<�<=D=�=�=�=k>�>?a?�?�?  �   0a0�0�0L1�1�12�2�2�2>3^3s3�3!4�4�4$5D5a5q5�5�5�5�5646d6�6�6�67$7D7a7�7�7�7808R8�8�8�8�89&9a9�9�9�9�9:�:�:�:�:�:�:;D;a;t;�;�;�;<D<d<�<�<�<�<�<'=b=�=�=�=2>`>�>�>�>�>!?4?d?�?�?�?�?     �   $0T0t0�0�01$1T1t1�1�1�1�1242F2a2t2�2�2�2�2�2343q3�3�3�3�3444T4q4�4�4�4�4�45$5D5d5�5�5�5�5616D6d6�6�6�6�67T7z7�7�7�78$8D8d8�8�8�8�89D9�9�9�9C:�:�:�:;D;q;�;�;�;�;<!<4<T<t<�<�<�<	==r=�=�=�=>$>D>�>�>�>�>�>?&?6?d?�?�?�?�?   0 �   000D0T0t0�0�0�0
1=1K1^1s1�1�1�1�1�12"222T2x2�2�2�2�2%3S3i3w3�3�3�3�3#494G4V4�4�4�4�4$5M5{5�5�5�56/6T6t6�6�6�6�67$7D7a7t7�7�7�7848T8t8�8�8�8�89!949Q9d9�9�9�9�9�9:%:6:H:a:4;b;�;�;<B<u<�<=E=U=�=�=1>m>�>�>5?r?�?�?   @ �   %0e0�0�051r1�1�12R2�2�23U3�3�34X4s4�4�4�4�455u5�5�556�6�67a7�7�7�7�788=8b8�8�8�8999x9�9�9:B:�:�:�:�:8;r;�;�;<�<�<�<�<=4=T=t=�=�=�=�=�=>>1>D>d>�>�>�>�>?$?A?d?�?�?�?�?   P �   040T0t0�0�0�01141T1q1�1�1�1�1242_2�2�2�2�233A3T3t3�3�3�3�3�344T4t4�4�4�4!5D5q5�5�5�5$6t6�67$7D7d7�7�7�7�7848D8t8�8�8�8949a9�9�9�9:1:T:�:�:�:;!;A;a;�;�;�;�;<!<A<a<�<�<�<�<=$=D=q=�=�=�=�=>2>T>q>�>�>�>�>?4?T?t?�?�?�?�?   ` �   $0D0d0�0�0�0�01A1�12D2t2�2�2�2313T3q3�3�3�3444d4�4�4�4.5r5�5�5�5�56D6q6�6�6�6�67D7t7�7�7�7848T8t8�8�8�8�89A9P9t9�94:a:t:�:�:�:;A;a;�;�;�;<!<A<d<�<�<�<$=T=�=�=�=>Z>�>�>�>?1?T?�?�?�?�?�? p �   0-0j0�0�01$1J1�1�12�23A3U3j3�3�3�34C4f4�4�4�4545x5�506t6�6�6�6797c7w7�7�7�78#8D8t8�8�8�89$9D9�9�9�9:1:Q:t:�:�:�:;T;�;�;�;<$<o<�<�<�<=.=X=s=�=�=�=>><>V>�>�>�>�>�>?O?c?x?�?�? � l   00A0[0{0�0�0g1z1�1�12212|2�4:7S7�7�7�7 878t8�8D:H:L:P:�:�:�:�:u;�;E<�<�<�<d=�=�=T>�>�>�>�>�>!?T? � $  �12a2h2�2�23:3I3t3}3�3�3�3�3�3�3�344(4F4e4w4�4�4�4�4�45"5/5G5Y5k5}5�5�5�5�5�56646F6X6a66�6�6�6�6�6$727?7W7i7{7�7�7�7�7�7�78(8D8V8h8q8�8�8�8�8�899-9N9d9�9�9�9�9�9�9::/:8:V:t:�:�:�:�:�:�:;;@;V;r;�;�;�;�;�;�;<<;<W<i<�<�<�<�<=1=�=�=�=�=�=�=> >1>:>M>�>�>�>?%?�?�?�?�?�? � �   -0O0d0�0�0�0�0�0�061H1�1�12q2�2�2�2�23A3T3t3�3�3�3�34t4b5i5p5w5~5�5�5�5�5�56�6E7�8�8�8k9�9�9�9::::!:(:/:6:=:D:K:R:Y:`:H;V;�;�;<w<�<�<�<�<�<X=x=�=�=�=�=d>�>�>�>�>?T?�?�?�?�?�?�?�? � �    0L0|0�0�0�0�01*1b1~1�1�1�1�1�1#2<2i2�2�2�23#3b3h3�3�3�3�3�3�34B4U4o4�4�4�4�4�4�4�5�5656{67E7�7�78V8�8�8"9X9�9�95:u:�:;E;�;�;"<R<�<�<�<%=u=�=�=>>:>b>�>�>5?�?�? � t   0e0�01U1�1�1"2b2�2�283�3�384�4�455�5�5%6u6�67X7�7X8�89U9�9�9%:u:�:;U;�;�;B<�<�<%=v=�=%>e>�>�>�>%?u?�?�? � @   E0�0�051�1�1F2�2�23U3�3�3%4u4�45E5�5�56D6�6�6?7�7<8   � 0   2<!<M<�<�<=U=�=�=>B>u>�>�>%?e?�?�?   � t   "0R0�0�0�01U1�1�152u2�2�253�3�3E4(6I6�8H9L9P9T9X9;:I:h:v:;;5;=;�;<0<><w<�<�=�=�=�=@>N>c>q>Q?d?�?�?�?�?     �   0D0c0v0�0�0�01A1T1�1�1�1�1$2d2�2�2�2�243T3q3�3�3�3�34D4v4�4�415D5t5�5�5�5�7�7�7 8�9�9:4:d:�:�:�:�:;$;T;�;�;�;�;�;<1<T<q<�<�<�<�=�=Z>_>�>�?�?�?  X   S0f0v0�0!1+1�1�1v2�2m3�334a4~4�4�46$6U6�6�6G7X7*;�;�;�<0=�=�=�=�=>>=>�>�>�?     �   0D0$1D1d1�1�12$2T2�2�2�2343�3�34$4+42494@4G4N4X4b4i4p4w4~4�4�4�4�4�4�4�4�4�45I5�5u699(979D9J9T9c9�9�9-:8:I:U:]:c:r:{:�:�:;;4;E;v;�;�;�;�;�;<'<;<�<�<�<�<�<�<�=�=%?2?E?e?o?�?�?�?�?�?   0 �   )090Q0r0�011.1>1J1]1d1o1u1�1�1f2373<3�5�5�56�6�6�6�67�8�9: :&:*:0:4:::>:D:H:M:S:W:]:a:g:k:q:u:�:�:�:;;';,;0;4;];�;�;�;�;�;�;�;�;�;�;<<<< <�<�<�<�<�<�<�<�<===D=H=L=P=T=X=\=`=�=�=�=�=�=P>d>�>?#?;?X?e?�?   @ `   S1e172A2N2i2p2�2�2�233g3m3~3�344*414�455.555�5�5�5�6�7�7�78W8�8�8�9M;�<>�>�>.?   P �   0u0z0�0�0�0�0�0$1*1E1u1�1�1�1)2�2�2�2w3�3�3�3�3�3n4�4�4�4�4-5>5�5�56666 6$6M6s6�6�6�6�6�6�6�6�6�6�67777v7�7�7�7�7�7�7�7�7-84888<8@8D8H8L8P8�8�8�8�8�8 99�9�9�9�9�9A:K:X:�:�:;;/;C;U;b;n;x;�;�;�;�;�<2=U=�=�>0?8?�?�? ` �   $000�0�0'131�1�1�1�2d4,5>5H5R5}5�5�5�5�5�5�5#6,686q6z6�6�6�6�6�7�7�7y8�8�8�8�8�8H9:7:�:�:;e;�;<<U<|<�<�<�<�<�<�<�<s=>l>�>�>�>?	?a?z?�?�?   p H   -0�0�1^2A4q4�4�45`5�5	6@6H6r78*8Z8d8p8y8�8g9_:t:;a=n=�=I>o?   � �   h0�0M2�3�6779:: :,:A:H:\:c:�:�:�:�:�:�:�:�:�:;;;#;);2;>;L;R;^;d;q;{;�;�;�;�;�;�;�;<[<a<�<�<�<�<�<e=�=�=�=�=>.>4>@>F>V>\>q>>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>
?????$?)?/?4?C?Y?d?i?t?y?�?�?�?�?�?�?�?�?�? � �   0a0l0�0�01111 1&1-141;1B1I1P1W1_1g1o1{1�1�1�1�1�1�1�1�1�1�1�1�1�1�12%2*2j3�3�315B5|5�5�5�5�5�5�5�5�56 636W6�6�6�6F7c7�7868�8�8�8�8�8�89979S9\9b9k9p99�9�9�9:1:T:g:�;j<�>c?�? � �   �4�5T7�7�7�7�7�7�7k9�9�9�9�9�9�9�9�9�9�9�9�9:	:::#:-:W:e:k:�:�:�:�:�:�:�:;�;�;�;�;>!>'>A>F>U>^>k>v>�>�>�>�>�>�>�>�>�>�>�>�>???&?-?3?A?H?M?V?c?i?�?�?�?�? � �   0�3�3�34K4�4c6n6v6�6�67�7�7�78k8}8�8�8�8�8�8�8�8�8�89(9:9H9]9g9�9�9�9�9�9+:�:;_;s;�;�;�;#<+<k<u<�<�<�<'=9=�=�=�=�=�=4?;?�?�?   � L   R01&12?2�2&45�5 66W6v67G7v7�78C8z8�89m9M:�:M<�<�<�<=@=o=n>�> � $   !0�0�0�0�01@1o1�2-3K3q3S:   � �   �4�4�455(5L5U5\5e5�5�5�5�56/6G6Y6}6�6�6�78#878@8m8�8�8�8�8�89'9:9E9J9Z9d9k9v99�9�9�9�9�9�9�93:@:j:o:z::�:);6;>;M;�;�;�;�;�;<<�=�=�=�=�=�=Y>_>u>�>�>�>�>�>�>=?P?�?�?�?�?�?�? � �   0�0�0�0�0|1�1�1�1�1�1�1�1 292A2N2�2�23$3?3K3W3c3�3�3�3�3�3�3�3�34
444(444=4F4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4@5�5�5�6�6'7-7d7�78�8�8�8�8�8�8�9`:;|;�;<<%<-<�<�<   X   �3	5$5u56 6B6}6�7�7-8�8�8�8�9�:�:�:�:;;%;B;n;�;�;�<�<�=�=�=>>>!>(>X>�>f?�?  t   ,0A0�0�0�0�0!1Y1�1�12!2E2h2�2�2�2�2�3�3�3�3�3�3�3-424w4|4�4�4�4�4555S;�;�;�;�;*<>=I=R=u=�=�=>>%>7>I>�>   L   �0�0�033-3J3y3�3�3�34\4�4�4)5N5�6:7�7�7>8G8�8�89$9=9�9�9�9�9?   @ �   G0K0O0S0W0[0_0c0g0k0o0s0w0{00�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�01�23/3N3�3�3�3�3*4:4g4o4�4�4�4�455)6�67)7�7�7�7i9�9?:^<m>v>�>�>x?}?�?�?�?�? P �   00Q0]0�0�0�0�01B1�2�3�3A4P4�4�4�5�5T6�6�6�6�7�7�78Q8�8N9{9�9�9�9�9�9�9�9�9
:::-:H:�:[;�;�;�;�;<'<B<b<�<�<= ={=�=�=�=�=>>>�>�>�>�>,? ` �   0)0/0?0D0\0b0q0w0�0�0�0�0�0�0�0�01,1I1�1�1�1�1�1�12!2)262=2�23r3	6o7�7�7�7�7)829�9�98:�:�<�<�<�<�<�<,=>�>�>�>H?[?v? p ,   �2�3;5j5�5r7n9r9v9z9~9�9�9�9�9�:�;)= � T   0�0 11/1A1T1f1�1�1�4�45,5I5T5k5�5�5\6�7�8]9S:[:;�;�<�<1=7=G=�=�=�>�?�?   � H   R041�1�1u2{2�2+3B3r3�3�6�61:5:9:=:A:E:I:M:Q:U:Y:]:j:D;^;m;�;�;< � 8   )6�7�7�7�7�7�788H9f9|:�:�:;a;�;�;�<�=�=�?�?   � L   030}0�0�0�1�1�1�1�1�1a2�2�23A3}3�3�3424�4K5�5�6q9�:�;�<?K?�?�?�? � h   @0�0�0I1�12T2�2]4�4i5�6!8t8�8�89B9s9�9�9&:v:�:�:�:I;�;�;�;)<c<�<�<�<*=_=�=�=�=*>Z>�>�>�>I?�?�? � P   0<0m0�0�0
1!1(1[1�1�1�1292\2�2�2�2�2333#3/393E3R3Z3d3v3�3�3�3�3�3�3 � �  `1d1h1l1p1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8�8�8�:�:�:�:�:�:�: ;;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======�=�=�=�=�=�>�>�>�> ??? � h    00P0T0X0\0`0d0h0l0|0�0�0@1D1H1L1P1T1X1\1t1x1|1P:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:,;0;4;8;�;�;     �   �9�9�9�9�9 :::: :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<  t  �2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 4444t6x677 7$7(707H7L7d7t7x7�7�7�7�7�7�7�7�7�7�7�788 8$8,8D8T8X8\8d8|8�8�8�8�8�8�8�8�8�8�8�8 999,90989P9`9d9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9 :::4:D:H:X:\:l:p:t:x:�:�:�:�:�:�:�:�:�:�:;;;;,;<;@;P;T;X;\;d;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�; << <0<4<D<H<L<T<l<|<�<�<�<�<�<�<�<�<�<�<�<�<�<===,=0=4=8=@=X=h=l=|=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>,>0>@>D>H>L>T>l>|>�>�>�>�>�>�>�>�>�>�>�> ???$?(?8?<?@?H?`?p?t?�?�?�?�?�?�?�?�?�?�?�?   �  0000 0$0,0D0T0X0`0x0�0�0�0�0�0�0�0�0�0�0�0�011 10141D1H1P1h1x1|1�1�1�1�1�1�1�1�1�1�1222 2$2,2D2T2X2h2l2t2�2�2�2�2�2�2�2�2�2�2�2 3333(383<3L3P3X3p3�3�3�3�3�3�3�3�3�3�3�3�3�3�344�5�5�5�5�56(6H6P6X6`6h6p6x6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7,747<7D7L7T7\7d7l7t7|7�7�7�7�7�7�7�7�7�78888$8,848<8D8P8p8x8�8�8�8�8�8�8�8�899(9H9P9\9|9�9�9�9�9�9�9�9:4:<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�:�:;$;,;4;<;D;L;T;\;h;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<d<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<====$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�> ???? ?(?0?8?@?H?P?X?`?h?p?x?�?�?�?�?�?�?�?�?�?�?�?�?�?   0 �  0000$0,040<0D0L0T0\0d0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1|1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2,242<2D2L2T2\2d2l2t2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3 4 4(444X4x4�4�4�4�4�4�4�4�4�4�4�4�4�4550585@5H5P5X5`5h5p5|5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6T6x6�6�6�6�6�6�6�6�6�6�677787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 8888 8(80888@8H8P8X8`8l8�8�8�8�8�8�8�8�8�8�8�8 9999 9,9L9T9\9d9l9t9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9::::$:,:4:<:H:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;d;�;�;�;�;�;�;�;�;�;�;�; <<<(<H<T<|<�<�<�<�<�<==,=@=H=`=l=�=�=�=�=�=�=>> >(>0><>\>d>l>t>|>�>�>�>�>�>�>???$?D?P?p?x?�?�?�?�?�?�?�?�?�?�?�? @ �  000040<0P0X0`0h0t0�0�0�0�0�0�0�0111 1@1D1H1P1d1l1�1�1�1�1�1�1�12$2P2X2|2�2�2�2�2�2�2�23,3<3P3`3t3|3�3�3�3�3�3�3 444<4L4`4h4�4�4�4�4�4�45$545@5`5p5|5�5�5�5�5�5606<6D6\6d6�6�6�6�6�6�67(707<7\7d7p7�7�7�7�7�7�7�7 888<8L8x8�8�8�8�8�8�8�8�89(949T9`9�9�9�9�9�9�9�9�9: :@:H:P:T:X:`:t:�:�:�:�:;;8;X;x;�;�;�;�;�;<8<X<d<p<�<�<�<�<�<�<�<== =P=X=\=t=x=�=�=�=�=�=�=�=�=�=�=>$><>@>\>`>�>�>�>�>�> ?? ?@?`?�?�?�?�?   P 0    0 0@0`0�0�0�0�0�0�0 1 1@1`1�1�1�1�1�1   ` 0   00 080<0@0\0x0�0�0�0�01L1�1�1�102P2�2�2 3 3@3d3�3�3�3�3�3�34 4<4h4l4p4t4�4�4�4�4�4�4�4�4�4�4�4 5555,5D5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6<6@6H6L6p6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6X7\7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7888@8x<�=�=�=>><>H>L>P>T>X>`>d>�?�?�?�?�?�?�?�?   p p   000181�3�34444$4,444<4D4L4T4\4d4l4t4|4�4�4�4�4�4�4N5R5V5Z5^5b5f5j5n5r5v5z5~5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�566
666666"6&6*6.62666:6>6B6F6J6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�677777 7$7(7,70747@7|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89999$9,949<9D9L9T9\9�9�9@:D:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        