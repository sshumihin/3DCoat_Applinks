MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       \��S�� �� �� ��h �� �k �� �} ��� ?,� �� �� x�� �z B�� �l �� �o �� Rich��                 PE  L {qP        � !	  ~  �      N,     �                         �                              �� S   � <                            0 �6  ��                            x� @            � \                          .text   �}     ~                   `.rdata  #^   �  `   �             @  @.data   �;   �     �             @  �.reloc  �B   0  D                 @  B                                                                                                                                                                                                                                                                                                                                                                                                U���V��H�QV�ҡ��H�U�AVR�Ѓ���^]� U���V��H�QV�ҡ��U�H�E�IRj�PV�у���^]� ����������U����P�E���   ��VWP�EP�E�P�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� ������������U��W�}��xS�]V�u����u��y�^[_]� ���������V���h� �N�����~ �N$�R\ ��^���������������V��N$����] �N��~ ��^�O� ���������������U���T  �\�3ŉE�Wj j�[ ����u_�M�3���� ��]�V������PWǅ����(  �x[ ����   ������Qj�h[ �����   ������RPǅ����$  �<[ ���}   ������P������h  Q�� ������h  R�� ���������P�I �@��u�+�$    ��/t��t������H��\uꍴ����V�U� h�V�� ����u.������PW�Z ���8���W� �^3�_�M�3���� ��]ËM�^3͸   _��� ��]���������3���������������3������������������������������j j j襦 �����U���\V��E�P�M�Q���E�   �E�    ��� �}� �  W�M��GZ ���B�P�M�Q�҃��E�Pj�M܍~Q������P�M��Z �U�R�M���] �M���Z ���H�A�U�R�Ћ��Q�J�E�P�у�h���M���Y �U�R�M���] �M��Z �E�j P�j �����M  ���Q�J�E�SP�ы��B�Pj j��M�h��Q�ҍE�P� ���Q�J�E�P�у�j ��蟃 ���B�P�M�Q�ҡ��H�Aj j��U�hx�R�ЍM�jQ�X �����B�P�M�Q���҃� j ����   hh��M������E�P�} ���Q�J�E�P���  h�h�   hh�   ���{� ����t	��轢  �3�WS�����  h�  ���Ԃ [�M��kY _^��]� j �U�R���E�   �E�    �h� [�M��?Y _^��]� �������U���SVW��j�~W�E�3�P�E�   �]��j� jW�M�Q���E�   �]��R� jW�U�R���E�   �]�蚍 jW�E�P���E�   �]��"� jW�M�Q���E�   �]��
� jW�U�R���E�   �]��� jW�E�P���E�   �]��ڌ jW�M�Q���E�   �]�� j
W�U�R���E�
   �]��
� j	�E�	   �]�W�E�P��蒌 jW�M�Q���E�   �]��z� jW�U�R���E�   �]��b� jW�E�P���E�   �]��J� jW�M�Q���E�   �]��2� _^[��]������������U���   V���� ��u^��]�SWh���M���V �E�P�M�Q�~$��j ��P�U�R��Z ��P���Z �M��gW �M��_W �M��WW 3ۉ^@��l SW�E���f ������  �E�P����W P�M��V jj�M�Q�M�htaoc��l ���M��E��W ���B�P�M�Q�҃�8]�t�E�P�nl ��_[3�^��]�Sh���M��������Q�R8�E�P�~j���ҡ��H�A�U�R�Ѓ��M��U �M�j	Q��j ��P�M��Y �M��pV h��M��U h���M��U �U�R�E�P�M�Q��l���R�Y ��P�E�P�Y ����l����#V �M��V �M��V �M�jQ�e ����t3�U�R�M��V ���QP�B8j���Ћ��Q�J�E�P���]Sh���M�����P�j ���B�P�M�Q�҃�Sh���M��W������P�R8�E�Pj���ҡ��H�A�U�R�Ћ��Q�B4��Sj���Ћ��Q�B0jj���Ћ��Q�B0jj���Ћ��Q�B0Sj���Ћ��Q�B0Sj���Ћ��Q�B0jj���Ћ��Q�B4Sj
���Ћ��Q�B0jj	���Ћ��Q�B0jj���Ћ��Q�B0Sj����Sh���M��]������Q�E�Pj�ϋR8�ҡ��H�A�U�R�Ћ��Q�B0��Sj���ЋM�W�p �M��j �M��GT �M��?T �M�Q�N$��T P�M��S �M�jj�U�Rhtaoc��i ���M��E��T ���H�A�U�R�Ѓ�8]�t�M�Q�ui ��_[3�^��]ËM�j�~W�{l �M��i ���E�   �]�B�P�M�Q�҃�SS�E�Pj�M�Q������P�U�R��襃 ���H�A�U�R�Ћ��Q�J�E�P�ы��E�   �]�B�P�M�Q�҃�SS�E�Pj�M�Q���0���P�U�R���D� ���H�A�U�R�Ћ��Q�J�E�P�у��E�   �]�h������B���   h  �Sjh���h  �Sj����P�E�P����} ��S�E�   �]�Q���   Sj����P�M�Q���� ��S�E�   �]�B���   Sj����P�E�P���� ��S�E�   �]�Q���   Sj����P�M�Q���T� ��S�E�   �]�B���   Sj����P�E�P���'� ���E�   �]�S�Q���   Sj����P�M�Q����� ��h���h  �Sjh���h  ��E�
   �]�B���   Sj
����P�E�P����| ��S�E�	   �]�Q���   Sj	����P�M�Q���� ��S�E�   �]�B���   Sj����P�E�P���]� ��S�E�   �]�Q���   Sj����P�M�Q���0� ���E�   �]�B�M̋PQ�҃�SS�E�Pj�M�Q�������P�U�R���� ���H�A�U�R�Ћ��Q�J�E�P�ы���S�E�   �]�B���   Sj����P�E�P���� h�  ����y �M�Q��e ��_[�   ^��]������������U���0V��~@ t~W�e �E��E�P�N$��P P�M��O jj�M�Q�M�htaoc��e �MЋ��P ���B�P�M�Q�҃���_t�������M���V�'l �M��e �E�P�Ve ��^��]���������������U���   SV��3�W�]��F@   �a����E����   ����   ���@  ���H�A�U�R�Ћ��Q�JSj��E�hh�P�эU�R�� ���H�A�U�R���	� h�h!  hh�   ����� ��,;�t���0�  ��VW���D�  _^�C[��]� ��3�VW���*�  _^�   [��]� �MQ�U�R���E�   �]��c� 9]�w  h�  ����w _^�   [��]� �k� h�h�   hj$���S� ��;�t�@   ��X�X�X�X�3���VW���O  ���H�A�U�R�Ћ��Q�JSj��E�h<�P�эU�R�� ���H�A�U�R�Ћ��Q�J�E�P�у� �U�Rj�E�P����������Q�J�E�P�ы��B���   ��Sj���҅�t1Sh���M��_������P�Rx�E�P�M��E�   ���E��u�]�E�t���H�A�U�R�Ѓ�8]�  �Q�������   ���Q�Bdj�M��Ћ��Q�����   h�Fh�   V�Ћ��Q��j���BhVW�M���j<��H���SQ�� ����H���RǅH���<   ��L�����P���ǅT���4���X�����`���ǅd���   ��h����T���uVSh��M��P����E�P�7 ���Q�J�E�P���(Sh��M��%����U�R� ���H�A�U�R�Ѓ����Q�J�E�P�у�_^�   [��]� �����U��V��N$����L �N��m ���=r �Et	V�� ����^]� ������������P�X����U�������M�P�P�P�P �P(�P0�P8�P@�PH�PP�XX���Q�P�Q�P�Q�P�Q�P�I�H�M��P�Q�P�Q�P �Q�P$�Q�P(�I�H,�M��P0�Q�P4�Q�P8�Q�P<�Q�P@�I�HD�M��PH�Q�PL�Q�PP�Q�PT�Q�PX�I�H\]� �����������U��M�U�A�
�E��B�I0���B�IH����A �
�A�A8�J���AP�J���X�A(�
�A�A@�J���AX�J���X�A�J�B �I0���B(�IH���X�A8�J �A �J���AP�J(���X �A@�J �A(�J���AX�J(���X(�A�J0�A0�J8���AH�J@���X0�A8�J8�A �J0���AP�J@���X8�A@�J8�A(�J0���AX�J@���X@�A�JH�BP�I0���BX�IH���XH�BP�I8�BH�I ���AP�JX���XP�A@�JP�BH�I(���AX�JX���XX]���U����UV��H�AVR�Ѓ���^]� ��������������U����H�U�I(��VWR�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]���U����E�H�U �E��VWR�UP�ERP�A$���U��$R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�,_��^��]��������������U���$�ESVW3ۍM�Q�M��]܉]�E�]��]��G$ �}S�U�R�E�P���, �M����: ;�th�����   �JX�E�P�ы���;�tJ�����   �PT���ҋ��Q|�M�RQPV�ҋ�����   ��U�R�Ѓ�_��^[��]� �����   �
�E�P�у�_^3�[��]� ������������U���$�EVW3��M�Q�M��}܉}�E�}��}��h# �MW�U�R�E�P�'+ �M����] ;�tZ�����   �JH�E�P�ы��u���B�HV�ы��B�HVW�ы����   ��M�Q�҃�_��^��]� ���H�u�QV�ҡ��H�QWj�h��V�ҡ����   ��U�R�Ѓ�_��^��]� ��������U���$�EVW3��M�Q�M��}܉}�E�}��}��x" �MW�U�R�E�P�7* �M����m ;�t8�����   �J8�E�P�ы������   ��M�Q�҃�_��^��]� �����   ��U�R�Ѓ�_3�^��]� �U���$�ESV3��u��M�Q�M��u܉u�E�u��u���! �MV�U�R�E�P�) ��t �����   �J�E�P�у���t��2ۍM�� ^��[t7�����   �P<�M�Q���]�����   ��U�R���E����]� �����   �
�E�P���E����]� ���������U���$�EVW3��M�Q�M��}܉}�E�}��}��! �MW�U�R�E�P��( �M����� ;�t[�����   �J@�E�P�ыu��H��P�N�H�V�P�@�N���V���   �
�F�E�P�у�_��^��]� ����u����   �V��^�M�Q�҃�_��^��]� U���$�EVW3��M�Q�M��}܉}�E�}��}��8  �MW�U�R�E�P��' �M����- ;�tD�����   �JL�E�P�ыu��P����C �����   ��M�Q�҃�_��^��]� �uW���JC �����   ��U�R�Ѓ�_��^��]� ����������U��Q���P�BdVWj�M�Ћ��Q�����   hX�Fh�  V�Ћ���j�E��QVP�Bh�M��N3���~S�]�I �M��R���AN G;�|�[�E�P�B� ���Q�J�EP�у�_^��]� �����U������H�AV�U�WR�Ћ��Q�Jj j��E�h��P�ы��B�Pd��j�M��ҋ���H���   hX�Fh�  V�ҋ���j�E��QVP�Bh�M���N3���~S�]���M��R���qM G;�|�[�E�P�r� ���Q�J�E�P�у�_^��]� �����U��Q�ESVW���   3�3�3�3ۃ��M�|#�@|�O���A�	�d$ p����u�E�M�;�}�@|��_�^�[��]� �����U����H�Q��   V�uV�ҡ��H�Qj j�hH�V�ҋE����
�  �$� / j hD��M��y����E�P���c  ���Q�J�E�P����  j h@���`����E�����`���R���gc  ��`����  j h8��M������M�Q���Bc  ���B�P�M�Q���p  j h4��M�������E�P���c  ���Q�J�E�P���?  j h0��M������U�R����b  �U��  j h(��M������M�Q���b  ���B�P�M�Q����   j h$��M��h����E�P���b  ���Q�J�E�P���   j h��M��7����U�R���\b  �U��   j h��M������M�Q���:b  ���B�P�M�Q���kj h���p����������p���P���b  ���Q�J��p���P���4j h���P���������P���R����a  ��P������H�AR�Ѓ����Q�J�E�P�ы��B�Pj j��M�h �Q�ҡ��P�B<�����Ћ��Q�RLj�j��M�QP���ҡ��H�A�U�R�Ѓ���^��]� �I �, �, - 5- f- �- �- �- . :. q. ����S�   V3�W���7�G�w�w�w�w�G(�w�w�w,�w$�w �G@�w0�w4�wD�w<�w8�GX�wH�wL�w\�wT�wP�Gp�w`�wd�wt�wl�wh���   �wx�w|���   ���   ���   �_���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   97t	W�(� ���7�w�w�w�w93t	S�� ���G0�3�s�s�s�s90t	P��� ���GH�w0�w4�wD�w<�w890t	P��� ���G`�wH�wL�w\�wT�wP90t	P�� ���Gx�w`�wd�wt�wl�wh90t	P�� �����   �wx�w|���   ���   ���   90t	P�g� �����   ���   ���   ���   ���   ���   90t	P�6� �����   ���   ���   ���   ���   ���   ��_^[����������SVW���� ���   3�93t	S��� ���3�s�s�s�s9��   ���   t	S�� ���3�s�s�s�s9wx�_xt	S�� ���3�s�s�s�s9w`�_`t	S�� ���3�s�s�s�s9wH�_Ht	S�b� ���3�s�s�s�s9w0�_0t	S�C� ���3�s�s�s�s9w�_t	S�$� ���3�s�s�s�s97t	W�	� ���7�w�w�w�w_^[�����U���  ��SVW���H�A�U�R�}��Ћ��Q�Jj j��E�hh�P�ы��B�P�M�Q�ҡ��H�Aj j��U�h\�R�ЋU��(�M�QR�E�P����P�M�Q�U�R��d  ��P�E�P��d  ���Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы]��S���B�H����V�ы��B�P�M�VQ�҃��������u�~ �E�    ��  3����H�A�U�R�Ћ��Q�Jj j��E�h��P�ы��B�P�M�Q�ҡ��H�Aj j��U�hX�R�Ћ��Q�J�E�P�ы��B�Pj j��M�hX�Q�ҡ��H�A��8���R�Ћ��Q�J��@j j���8���hT�P�ыF���D8��j0j jǋB�P$j ���������$Q�ҋء��H������AR�Ћ��Q�J�����PS�ы��B�P������Q�ҋF�D8��,j0j ǡ��H�A$jj ���������$R�Ћ��Q�J�؍�(���P�ы��B�P��(���QS�ҡ��H�A������R�ЋF���8�Q�J$��,j0j j�j ��������$P�ы��؋B�P��H���Q�ҡ��H�A��H���RS�Ћ��Q�J�����P�ы��B�P�M�Q�ҡ��H�I�U�R��8���P�ы��B�P<��8�M��ҋ��Q�RLj�j���H���QP�M��ҡ��H�A�U�R�Ћ��Q�R�E�P�M�Q�ҡ��P�B<���M��Ћ��Q�RLj�j��M�QP�M��ҡ��H�A��h���R�Ћ��Q�R��h���P�M�Q�ҡ��P�B<����h����Ћ��Q�RLj�j���(���QP��h����ҡ��H�A�U�R�Ћ��Q�R�E�P��h���Q�ҡ��P�B<���M��Ћ��Q�RLj�j��M�QP�M��ҡ��H�A��x���R�Ћ��Q�R��x���P�M�Q�ҡ��P�B<����x����Ћ��Q�RLj�j������QP��x����ҡ��H�A��X���R�Ћ��Q�R��X���P��x���Q�ҡ��P�B<����X����Ћ��Q�RLj�j��M�QP��X����ҡ��H�I�U�R��X���P�ы��B�P��X���Q�ҡ��H�A��x���R�Ћ��Q�J�E�P�ы��B�P��h���Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P��H���Q�ҡ��H�A��(���R�Ћ��Q�J�����P�ы��B�P��8���Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҋE���Q��<P�B����S�Ћ��Q�J�E�SP�ыM܃������E�@��;F�E��j����}܋]���B�P�M�Q�ҡ��H�Aj j��U�hh�R�Ћ��Q�J�E�P�ы��B�Pj j��M�hL�Q�ҡ��H�U�I(R�����P�ы����B�P�M�Q�ҡ��H�A�U�RV�Ћ��Q�J�����P�ы��B�P�M���@Q�ҡ��H�I�U�R�E�P�ы��B�P<���M��ҋ��Q�RLj�j��M�QP�M��ҡ��H�A�U�R�Ћ��Q�R�E�P�M�Q�ҡ��P�B<���M��Ћ��Q�RLj�j��M�QP�M��ҡ��H�I�U�R�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ���S����Q�BV�Ћ��Q�J�E�VP�у����m���S���������B�P�M�Q�҃�_^[��]� �������U���  ��SVW���H�A�U�R�}��Ћ��Q�Jj j��E�h��P�ы��B�P�M�Q�ҡ��H�Aj j��U�h\�R�Ћu�F,��(�M�QP�U�R����P�E�P�M�Q��[  ��P�U�R��[  ���H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�ЋM�����BQ�H����S�ы��B�P�M�SQ�҃����'���3�9]�]��  ���H�A��(���R�Ћ��Q�Jj j���(���h��P�ы��B�P������Q�ҡ��H�Aj j�������hX�R�Ћ��Q�J������P�ы��B�Pj j�������hX�Q�ҡ��H�A��h���R�Ћ��Q�J��@j j���h���h��P�ыF����j0�<[�j �j��D8ǋB�P$j ���������$Q�҉E����H�A������R�Ћ��Q�M��R������PQ�ҡ��H�A������R����F�d8���Q�J$��,j0j �jj ���������$P�ы��E��B�P������Q�ҡ��H�E��I������RP�ы��B�P������Q�ҋF�8��,j0j ǡ��H�A$jj ���������$R�Ћ��Q�J�E���H���P�ы��B�U��@��H���QR�Ћ��Q�J������P�ы��B�P��8���Q�ҡ��H�I��8���R��h���P�ы��B�P<��8��8����ҋ��Q�RLj�j���H���QP��8����ҡ��H�A��X���R�Ћ��Q�R��X���P��8���Q�ҡ��P�B<����X����Ћ��Q�RLj�j�������QP��X����ҡ��H�A��x���R�Ћ��Q�R��x���P��X���Q�ҡ��P�B<����x����Ћ��Q�RLj�j�������QP��x����ҡ��H�A������R�Ћ��Q�R������P��x���Q�ҡ��P�B<���������Ћ��Q�RLj�j�������QP�������ҡ��H�A������R�Ћ��Q�R������P������Q�ҡ��P�B<���������Ћ��Qj�j�������QP�RL�������ҡ��H�A������R�Ћ��Q�R������P������Q�ҡ��P�B<���������Ћ��Q�RLj�j���(���QP�������ҡ��H�I�U�R������P�ы��B�P������Q�ҡ��H�A������R�Ћ��Q�J������P�ы��B�P��x���Q�ҡ��H�A��X���R�Ћ��Q�J��8���P�ы��B��H���Q�P�ҡ��H�A������R�Ћ��Q�J������P�ы��B�P��h���Q�ҡ��H�A������R�Ћ��Q�J������P�ы��B�P��(���Q�ҋE���Q��<P���ĉE�P�B�Ћ��Q�E��RP�M�Q�ҋM����������H�A��x���R�Ћ��Q�Jj j���x���h��P�ы��B�P������Q�ҡ��H�Aj j�������hX�R�Ћ��Q�J������P�ы��B�Pj j�������hX�Q�ҡ��H�A�����R�Ћ��Q�J��@j j������h��P�ыV�D:(��j0j �D:���H�A$jj ����X����$R�Ћ��Q�J�E�������P�ы��B�U��@������QR�Ћ��Q�J��X���P����V��,�D:�`���H�A$j0j jj ��������$R�Ћ��Q�J�E���8���P�ы��B�U��@��8���QR�Ћ��Q�J�����P�ыV���D:�H�A$��,j0j j�|:j ����8����$R�Ћ��Q�J��������P�ы��B�P������QW�ҡ��H�A��8���R�Ћ��Q�J�E�P�ы��B�M�Q������@R�Ћ��Q�B<��8�M��Ћ��Q�RLj�j�������QP�M��ҡ��H�A��(���R�Ћ��Q�R��(���P�M�Q�ҡ��P�B<����(����Ћ��Q�RLj�j�������QP��(����ҡ��H�A��H���R�Ћ��Q�R��H���P��(���Q�ҡ��P�B<����H����Ћ��Q�RLj�j���8���QP��H����ҡ��H�A��H���R�Ћ��Q�R��H���P��H���Q�ҡ��P�B<����H����Ћ��Q�RLj�j�������QP��H����ҡ��H�A������R�Ћ��Q�R������P��H���Q�ҡ��P�B<���������Ћ��Q�RLj�j�������QP�������ҡ��H�A��h���R�Ћ��Q�R��h���P������Q�ҡ��P�B<����h����Ћ��Qj��RLj���x���QP��h����ҡ��H�I�U�R��h���P�ы��B�P��h���Q�ҡ��H�A������R�Ћ��Q�J��H���P�ы��B�P��H���Q�ҡ��H�A��(���R�Ћ��Q�J�E�P�ы��B�P������Q�ҡ��H�A��8���R�Ћ��Q�J������P�ы��B�P�����Q�ҡ��H�A������R�Ћ��Q�J������P�ы��B�P��x���Q�ҋE���Q��<P�B����W�Ћ��Q�J�E�WP�ыM����C������B�P�����Q�ҡ��H�Aj j������h��R�Ћ��Q�J������P�ы��B�Pj j�������hX�Q�ҡ��H�A��(���R�Ћ��Q�Jj j���(���hX�P�ы��B������Q�P�ҡ��H�A��@j j�������h��R�ЋF���Q�J$��j0�|[�j �j��D8�j ����x����$P�ы��E��B�P������Q�ҡ��H�E��I������RP�ы��B�P��x���Q����F�d8��,j0j ǡ��H�A$jj ����h����$R�Ћ��Q�J�E���X���P�ы��B��X���Q�U��@R�Ћ��Q�J��h���P�ыF���8��,j0j jǋB�P$j ����H����$Q�ҋ����H�A������R�Ћ��Q�J������PW�ы��B�P��H���Q�ҡ��H�A��X���R�Ћ��Q�R��X���P������Q�ҡ��P�B<��8��X����Ћ��Q�RLj�j�������QP��X����ҡ��H�A��x���R�Ћ��Q�R��x���P��X���Q�ҡ��P�B<����x����Ћ��Q�RLj�j���(���QP��x����ҡ��H�A������R�Ћ��Q�R������P��x���Q�ҡ��P�B<���������Ћ��Q�RLj�j���X���QP�������ҡ��H�A������R�Ћ��Q�R������P������Q�ҡ��P�B<���������Ћ��Qj�j�������Q�RLP�������ҡ��H�A��h���R�Ћ��Q�R��h���P������Q�ҡ��P�B<����h����Ћ��Q�RLj�j�������QP��h����ҡ��H�A�����R�Ћ��Q�R�����P��h���Q�ҡ��P�B<��������Ћ��Q�RLj�j������QP������ҡ��H�I�U�R�����P�ы��B�P�����Q�ҡ��H��h����AR�Ћ��Q�J������P�ы��B�P������Q�ҡ��H�A��x���R�Ћ��Q�J��X���P�ы��B�P������Q�ҡ��H�A��X���R�Ћ��Q�J������P�ы��B�P������Q�ҡ��H�A��(���R�Ћ��Q�J������P�ы��B�P�����Q�ҋE���Q��<P�B����W�Ћ��Q�J�E�WP�ыM����R����V|�E�<���  ���H�A�U�R�Ћ��Q�Jj j��E�h��P�ы��B�P�M�Q�ҡ��H�Aj j��U�hX�R�Ћ��Q�J�E�P�ы��B�Pj j��M�hX�Q�ҡ��H�A������R�Ћ��Q�J��@j j�������h��P�ыF����j0�|[	�j �j��D8ǋB�P$j ����(����$Q�҉E����H�A������R�Ћ��Q�M��R������PQ�ҡ��H�A��(���R����F�d8���Q�J$��,j0j �jj ��������$P�ы��E��B�P�����Q�ҡ��H�E��I�����RP�ы��B�P�����Q�ҋF�8��,j0j ǡ��H�A$jj ���������$R�Ћ��Q�J�������P�ы��B�P�����QW�ҡ��H�A������R�Ћ��Q�J�E�P�ы��B�@�M�Q������R�Ћ��Q�B<��8�M��Ћ��Q�RLj�j������QP�M��ҡ��H�A�U�R�Ћ��Q�R�E�P�M�Q�ҡ��P�B<���M��Ћ��Q�RLj�j��M�QP�M��ҡ��H�A������R�Ћ��Q�R������P�M�Q�ҡ��P�B<���������Ћ��Q�RLj�j������QP�������ҡ��H�A������R�Ћ��Q�R������P������Q�ҡ��P�B<���������Ћ��Q�RLj�j��M�QP�������ҡ��H�A�����R�Ћ��Q�R�����P������Q�ҡ��P�B<��������Ћ��Qj�j�������QP������RL�ҡ��H�A��8���R�Ћ��Q�R��8���P�����Q�ҡ��P�B<����8����Ћ��Q�RLj�j��M�QP��8����ҡ��H�I�U�R��8���P�ы��B�P��8���Q�ҡ��H�A�����R�Ћ��Q�J������P�ы��B�P������Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P�����Q�ҡ��H�A�����R�Ћ��Q�J������P�ы��B�P������Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҋE���Q��<P�B����W�Ћ��Q�J�E�WP�ыM��������E�V|�@;E�E�j����}����H�A�U�R�Ћ��Q�Jj j��E�h��P�ы��B�P�M�Q�ҡ��H�Aj j��U�hL�R�Ћ��v,�Q�J(������VP�ы����B�P�M�Q�ҡ��H�A�U�RV�Ћ��Q�J������P�ы��B�P�M؃�@Q�ҡ��H�I�U�R�E�P�ы��B�P<���M��ҋ��Q�RLj�j��M�QP�M��ҡ��H�A�U�R�Ћ��Q�R�E�P�M�Q�ҡ��P�B<���M��Ћ��Q�RLj�j��M�QP�M��ҡ��H�I�U�R�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ]��S������Q�BV�Ћ��Q�J�E�VP�у�������S���������B�P�M�Q�҃�_^[��]� �������������U���  ���USVWj ��HH��p  h�  R�Ћ��Q�}��j �E����   j���Ћ��Qj �E����   j���Ћ��Q�J���E�P�}��у�����  �~ ��  ��h���� �����R�j� ��胯 P��h���� ������l ���H�A�U�R�Ћ��Q�Jj j��E�h��P�у��U�R��h����� ���H�A�U�R�Ћ��Q�J�E�P�ы��B�Pj j��M�h��Q�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h��P�у�,�U�R�E�P�����Q��h����g ���` P�U�R�E�P��?  ��P�M�Q��?  ���J�U�RP�A�Ћ��Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ѓ� ������/ ���Q�J�E�P�ы��B�P�M�Q�ҋ]���H�Q��S����W�ҡ��H�A�U�WR�Ѓ��������S��������h����� ��]���Q�J�E�P�ы��B�Pj j��M�h��Q�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h��P�ы����   �M�Px��(�ҍM�QP�U�R�E�P�>  ��P�M�Q�>  ���J�U�RP�A�Ћ��Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�у�$���B�HS����W�ы��B�P�M�WQ�҃�������S���W����E�}PWS���w����}� t�M��UQRWS���P������H�A�U�R�Ћ��Q�Jj j��E�h��P�ы��B�P�M�Q�ҡ��H�Aj j��U�h\�R�ЋU��(�M�QR�E�P�t���P�M�Q�U�R�V=  ��P�E�P�I=  ���Q�R�M�QP�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��J�Q��(S����P�E�ҡ��H�U�IR�E�P�у����d������B�P��X���Q�E    �ҡ��H�Aj j���X���h��R�Ћ��Q�J�E�P�ы��B�Pj j��M�h��Q�҃�(�} �E    �U  �}� ��  �~ ��  ���   �M�������   ����� ���   �ȋBx�Ћ��Q�R�M�QP�ҡ��P�Rx����X���P�M��҅��8  ���H�A�U�R�Ћ��Q�Jj j��E�h��P�ы��B�P�M�Q�ҡ��H�Aj j��U�h��R�Ѓ�(�M�Q�U�R�E�P������Q�A;  ��P������R�1;  ���Q�R�M�QP�ҡ��H�A������R�Ћ��Q�J������P�ы��B�P�M�Q�ҡ��H�A�U�R�Ѓ�$S���ĉE���QP�B�Ћ��Q�E�RP�M�Q�҃����W������H�I��X���R�E�P�у����B�P��H���Q�ҡ��H�Aj j���H���h��R�Ћ��Q�R�E�P��H���Q�ҡ��H�A��H���R�ЋO|�U�� �<� �E    �o  �]�ۡ��H�A��8���R�Ћ��Q�Jj j���8���hX�P�ы��B�P<���M��ҋ��Q�RLj�j���8���QP�M��ҡ��H�A��8���R�ЋG4��VÍD���Q�J(P�����P�ы��E�B�P��(���Q�ҡ��H�E�I��(���RP�ы��B�P�����Q�ҡ��P�B<���M��Ћ��Qj�j���(����RLQP�M��ҡ��H�A��(���R�Ѓ��}� �  �\ �  ���Q�J�E�P�ы��B�Pj j��M�h��Q�ҡ��P�B<���M��Ћ��Q�RLj�j��M�QP�M��ҡ��H�A�U�R�ЋGL��NÍD���Q�J(P��t���P�ы��E�B�P�M�Q�ҡ��H�E�I�U�RP�ы��B�P��t���Q�ҡ��P�B<���M��Ћ��Qj�j��M��RLQP�M��ҡ��H�A�U�R�Ѓ��E�O|�U@��;��E������]���H�A�U�R�Ћ��Q�Jj j��E�h��P�ы��B�P<���M��ҋ��Q�RLj�j��M�QP�M��ҡ��H�A�U�R�Ћ��Q��S���ĉEP�B�Ћ��Q�E�RP�M�Q�҃��������E�O|��U@;E�E��������H�A�U�R�Ћ��Q�Jj j��E�h��P�ы��B�P�M�Q�ҡ��H�Aj j��U�hL�R�Ћ��Q�E�R(P��t���Q�ҋ����H�A�U�R�Ћ��Q�J�E�PW�ы��B�P��t���Q�ҡ��H�A�U���@R�Ћ��Q�R�E�P�M�Q�ҡ��P�B<���M��Ћ��Q�RLj�j��M�QP�M��ҡ��H�A�U�R�Ћ��Q�R�E�P�M�Q�ҡ��P�B<���M��Ћ��Q�RLj�j��M�QP�M��ҡ��H�I�U�R�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ���S�����Q�BW�Ћ��Q�J�E�WP�у�������S���4������B�P�M�Q�ҡ��H�A��X���R�Ћ��Q�J�E�P�у�_^[��]� U�����   SV��H�A�U�WR�Ћ��Q�Jj j��E�hX�P�ы��B�P�M�Q�ҡ��H�I�U�R�EP�ы��B�P<�� �M��ҋ��Q�RLj�j��M�QP�M��ҡ��H�A�U�R�ЋM�]��QS�U�R���
������H�A�U�R�Ћ��Q�Jj j��E�h��P�ы��B�P�M�Q�ҡ��H�Aj j��U�hX�R�Ћ��Q�J�E�P�ы��B�Pj j��M�hX�Q���E���<�E�Pj0j jj ���M��$Q�����E���P�U�Rj0j jj ����x����$P�����E���P�M�Qj0j jj ����\����$R�Z�����P�� ���P��2  ��P�� ���Q��2  ��P��@���R�2  ��P�����P�2  ��P��0���Q�2  �����B�P<���M��ҋ��Qj�j�WP�BL�M��Ћ��Q�J��0���P�ы��B�P�����Q�ҡ��H�A��@���R�Ћ��Q�J�� ���P�ы��B�P�� ���Q�ҡ��H�A��\���R�Ћ��Q�J��x���P�ы��B�P�M�Q�ҡ��H�UЋAR�Ћ��Q�J�E�P�ы��B�P�M�Q�ҋE���Q��,P�B����W�Ћ��Q�J�E�WP�у��������Uh�  RS���<������4  h�  P��P���P���0����M��� �M�Q��l����� �MP��P���R�E�P�e� P菿 ���M�� ��l���� ���Q�J�E�P�ы��B�Pj j��M�hX�Q�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h��P�у�(�U�R�EP�M�Q��x���R�u0  ��P�E�P�h0  ���Q�R�M�QP�ҡ��H�U��AR�Ћ��Q�J��x���P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ы��B�Pj j��M�h��Q�҃�8�E�P��x���Q�M��) P�U�R�/  �����P�B<���M��Ћ��Qj�j�WP�BL�M��Ћ��Q�J�E�P�ы��B�P��x���Q�ҡ��H�A�U�R�ЋM���B��Q�H����W�ы��B�P�M�WQ�҃���������M�� ��P���� ���H�A�U�R�Ћ��Q�J�EP�у�_^[��]�$ �U����   SV��W�M��z ���H�A�U�R�Ѓ��M�Q�Mj�U�R�D���P��8���� ��8���P�M�� ��8���� ���Q�J�E�P�ы��B�P�M�Q�ҋM���E�P�� P�M��� �M��� ���Q�J�E�P�ы��B�P3�Sj��M�h��Q�҃��E�P�M��M ���Q�J�E�P�у��U�R�M��< P�&� ���H�A�U�R�Ѓ��-	 h1D4ChCD4C�E����ɸ PSj�M�Q���J	 ��u"�U�R�	 ���M��]�� 3�_^[��]� �F;É]�  �F�M���<��B�P�M�Q�ҡ��H�A��t���R�Ћ��Q�Jj j���t���h��P�ы��B�P��T���Q�ҡ��H�Aj j���T���h�R�Ћ����   �Bx��,���Ћ��Q�J�؍E�P�ы��B�@�M�Q��T���R�Ћ��Q�B<���M��Ћ��Qj�j�SP�BL�M��Ћ��Q�J�E�P�ы��B�@�M�Q�U�R�Ћ��Q�B<���M��Ћ��Q�RLj�j���t���QP�M��ҡ��H�I�U�R�E�P�ы��B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J��T���P�ы��B�P��t���Q�ҋE����Q��P�B����S�Ћ��Q�J�E�SP�у����F������B�P��d���Q�ҡ��H�Aj j���d���h��R�Ћ��Q�R�E�P��d���Q�ҡ��H�A��d���R�ЋM����B�� Q�H����S�ы��B�P�M�SQ�҃���诽��h�  W��袺����tG���H�Q����S�ҡ��H�Qj j�h��S�ҋE��M��h4  h@  WPQ������h�  W���J�����tI���B�H����S�ы��B�Hj j�h��S�ыU��E��h�	  hD  WRP���������Q�J��D���P�ы��B�Pj j���D���h�Q�ҡ��H�I�U�R��D���P�ы��B�P��D���Q�ҋE����Q�� P�B����W�Ћ��Q�J�E�WP�у����e������B�P�M�Q�ҡ��H�Aj j��U�hԔR�Ћ��Q�R�E�P�M�Q�ҡ��H�A�U�R�ЋM��� Q���B�H����W�ы��B�P�M�WQ�҃����ڻ�����H�A�U�R�Ћ��Q�Jj j��E�hȔP�ы��B�@�M�Q�U�R�Ћ��Q�J�E�P�ыU����H�� R�Q����W�ҡ��H�A�U�WR�Ѓ����P����M�Q���������B�P�M�Q�ҋE@��;F�E������M��( �E�P�� ���M��E�    ���  _^�   [��]� ���������������U���  SVW��hG  �]��� �K 3����������;���  ��������  ���H�A�U�R�Ћ}���M�Qj�U�R���Z���P�M����  �E�P�������2 �M��:�  ���Q�J�E�P�ы��B�P�M�Q�ҋM���E�P�� P������� �M����  ���Q�J�� ���P�ы��B�PVj��� ���hp�Q�҃��� ���P�������\  ���Q�J�� ���P�у���l�����  ���B�M�Q�P�҃��E�Pj�M�Q���c���P�M����  �U�R��l����;  �M��C�  ���H�A�U�R�Ћ��Q�J�E�P�у�hd��M��P�  �U�R��l����  �M����  ���������  ���H�A�U�R�Ѓ��M�Qj�U�R���ɞ��P�M��@�  �E�P��������  �M���  ���Q�J�E�P�ы��B�P�M�Q�҃�hX��M���  �E�P�������v�  �M��^�  �M�Q��������  P��� ���B�P�M�Q�҃��E�P��l������  P�ϱ ���Q�J�E�P�у��U�R��������  P襱 ���H�A�U�R�����U����U��M��P�Q�]��U�R��x����U�P�荍�����U�Qݝx����������U�ݕ����ݕ����ݕ����ݕ����ݝ����谯�������   ���   �ыMVP�E�诏 �����   �M􋐐   �҅��%  �  h1D4ChCD4C�E��E�覯 �M�PVj������P�#  ��uV�M�Q���  ���u����   ���   �M�Q�҃��u􍍈������  ��l������  ���������  3�_^[��]� Vh���M��k����E�P����M�Q�U�R�������O�  PV��#  ����螶�����H�A�U�R�Ћ��Q�J�E�P�у�j h���M��	����U�R����E�P�M�Q��l������  PV�#  �����<������B�P�M�Q�ҡ��H�A�U�R�Ѓ�j h���M�觛�����Q���   �u�j j����V����M�QP�U�R��觷��PV�#  �����Ƶ�����H�A�U�R�Ћ��Q�J�E�P�ы��B���   ��3�Vj����;�t�E�P����Vh@��������i������Q���   Vj����;�t�M�Q����Vh0��ۚ�����4������B���   Vj����P�E�P������P蜮 ���Q�J�E�P�ыM������  Vh ��M�聚��Vh��M��s����U�R�����P�������]�  P�M�Q������R��!  ��P������P��!  P�&� ���Q�J������P�ы��B�P������Q�ҡ��H�A�����R�Ћ��Q�J�E�P�ы��B�P�M�Q�҃�$���  h1D4ChCD4C�E��E��w� �M�PVj������P���  ��u(�M�Q��  �U�R�u���  ���M�u��M  ��������H�A�� ���R�Ѓ�Vh���M��S������Q�R�� ���P�M�Q�ҡ��H�A�U�R�ЋM���Q���� �����R�������j����   �E��E��E�P�E��  �u��u��u��� ��Vh���M��՘��Vh��M��ǘ���M�Q�U�R�����hЕP�� P�M�Q������R�=   ��P������P�-   ��P�� �����������Q������P�J�ы��B�P������Q�ҡ��H�A�����R�Ћ��Q�J�E�P�ы��B�P�M�Q�ҋE���P���� �����R�ԗ�����]���Vh���M�����Vh���M�������� �M�QP�����R�y���P�E�P������Q�X  ��P������R�H  ��P�� ����������H�A������R�Ћ��Q�J������P�ы��B�P�����Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�ыU���R���� �����P�������y����M�Q���������B���   Vj���ҋM�s�s�Eġ����   ���   �u��Ѕ��c  虫 �����   �E��M􋒔   P�ҋ�����   �B�Ήu���=�  ��  ���Q�J������P�ы��B�Pj j�������h��Q�ҡ����   �Bx������P������Q������R��  P�*� ���H�A������R�Ћ��Q�J������P�у��������������B�P������Q�ҡ��H�Aj j�������h��R�Ћ����   �Bx������P������Q������R�7  P聩 ���H�A������R�Ћ��Q�J������P�у��}� ��  ���BH���   h�  V�у�P��<����5  j��T����(  j ��<����K  ���E�    �-� ���}ȅ���  �����   �P����=�  ��  hF  h�  W���`������i  j ���E�   ��� ������  h�  W�E�P���������Q�B<�M��Ѕ���   V��T����  �M��� ������   ��    �����   �B����=)  ��   �����   �Bx���Ћ��Q�Rx�M�Q���҅�ui���� �؍E�P������Qh���3�V���D� ��tB������F;E��d$ ��h�����@���J��@;E�~�U�R������Ph���V���� ��u������   �B(���Ћ����1������X����1j ��<����  ���B�P�M�Q�ҋ]��}ȃ������   �B(���Ћ��Eȅ��@�����X����9 ��   ���B�P�M�Q�ҡ��H�Aj j��U�h��R�Ћ����   ��������@|���U�R�Ћ��Q�J�E�P�ы���JT�Q3�WP�҃�;���  �����Q���&� ����U��U��M��]�Q�B�PHh�  ������ҋ�X����������� �}� ��   ��h��� �E�    ��   3�9s~X�d$ �S����� ���   �ȋBx�Ћ�X����U����������   �Bx�Ћ��Q�ȋBxW�Ѕ�t1F;s|��s��X����U��<���|jjjV���+  ��t�C�<��E�@;�h����E��c������QH�u܋�p  j h�  V�Ћ��QHj ��������p  h�  V�Ћ��QH���������   h�  V�Ћ��QH�����   h�  V�}��Ћ���4�����(�u�;�t(}+�PV�� ����w  �jj��+�QP�� ����`  3���~9����������������3�;Q��$�����@����;Eȉ\��������|ԋ}�������P��胬����8���������;�t ������}+�PW��  �jj+�WP��  ���QH�M܋R8��X���P�ҋ�   �����������P������Q��$���R肣����݅|���3ۃ}�݅t���݅l���݅d���݅\���݅T����  �}�����������B(����G��    ݅<����������H؍t��܅$������H������H����]�݅D����H�܅,������H������H����]�݅L����H�܅4������H������H����E���E��Y�Y������݅<����L1�H�܅$������H���������]�݅D����H�܅,������H���������]�݅L����H�܅4������H���������E���E��Y�Y݅<����H܅$������H�����H���������L��]�݅D����H܅,������H�����H���]�݅L����H܅4������H�����H���E���E��Y�Y������݅<����L �H ȃ�`��܅$������H������H���ݝ����݅D����H�܅,������H������H���ݝ���݅L����H�܅4������H������H���݅�����]�݅������]��E���Y�E��Y����;]���   �������[�D��U�����+�+�݅<����������H��ȃ���܅$������H������H���ݝ����݅D����H�܅,������H������H���ݝ���݅L����H�܅4������H������H���݅�����]�݅������]��E���Y�E��Y�e�����8����݋���������������;�t&}+�QP�������l  �jj+�PQ�������W  �]�3�3Ʌ���   ��������$��������$    �<�������u.�r�4��2�������t��r��������t��r��������t���2�4��r��������t��r��������t���$����A��;�|����B�M���   j j�҅��X  ���HH�u܋��   j h'  V�ҋ������Y  ��8���������;�t,}+�QP�������]  �jj+�PQ�������X  ��8��������;�t&}+�QP�������'
  �jj+�PQ�������  ���k� ��ݕ$���3�ݕ,���3�ݕ4���������ݕ<���ݕD���ݕL���ݕT���ݕ\���ݕd���ݕl���ݕt���ݝ|������a  ���HD�������I,��$���RWP�ы�$����v�Ƀ�Ƀ<��7  ��������l������p����T��t����T��x����T��|����T�U��T��������D��T������X����P��\����H��`����P��d����H��h����P�������N�I��<������@����P��D����P��H����P��L����P��P����P�������V�R�Ë�$������(����X��,����X��0����X��4����X��8����X�������4��������F�D��������]ȉ�����������   �������
��T������X����P��\����P��`����P��d����P��h����P�������D��<������@����P��D����H��H����P��L����H��P����P�������N�I��$������(����P��,����P��0����P��4����P��8����P�������4��������V�T�����������$���4�G;�������M��E��}�u�SQ�M܍�����RPQW�������������V���P���   j j���Ѕ�t	������N������赩���ދ��u����   �M􋐐   F�u���;������3��M����  9u�t9s~�EWP���������Q�J�� ���P�эU�R�O�  �E�P�u��C�  ���  j h���������	���3�Vh|��M�����������   �M܋Bx�Ѝ�����QP�U�R������P�n  ��P������Q�^  P訛 ���B�P������Q�ҡ��H�A������R�Ћ��Q�J�E�P�ы��B�P������Q�҃� �������z������H�A�� ���R�ЍM�Q�]�  �U�R�u��Q�  ���M�u���  �y����������3������H�A�� ���R�ЍM�Q��  �U�R�}��
�  ���}����   ���   �U�R�Ѓ��}�� ������Q�J�E�P�ы��B�P3�Wj��M�hH�Q�ҡ��H�A�U�R�Ћ��Q�JWj��E�h<�P�ы����   �Px��(���ҋ���H�A������R�Ћ��Q�R������P�M�Q�ҡ��P�B<���������Ћ��Qj�j�VP�BL�������Ћ��Q�J�����P�ы��B�@�����Q������R�Ћ��Q�B<��������Ћ��Q�RLj�j��M�QP������ҍ����P�v� ���Q�J�����P�ы��B�P������Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�у��������K������B�P�� ���Q�ҍE�P�-�  �M�Q�}��!�  ���}����   ���   �M�Q�҃��}��6������Q�J�E�P�ы��B�PVj��M�h$�Q�ҍE�P薘 ���Q�J�E�P�у�������R�5� �����   ���   �U�R�Ѓ��������u���  ��l�����  ��������  _^�   [��]� ��������̡�V�񋈈   ���   V�҃��    ^���������������VW��3�9>t	V�k ���>�~�~�~�~_^�������������U��Q3�9A~V�u�2@��;A|�^]� ���������������U��EV���
�   ^]� �MW��|/�~;�}(�> t#�~ u%���H��0  h��h�  �҃�_3�^]� ��;�|���;���_�   ^]� S�;�|�ߋ�+���;ȉ]��   ^��~�F�I���QP�[��P�d� ���N��~;ύI�ЉV�'  ������V+ӍR���R��)F+ȍ@��N�N�Q�+�Q�� �F���Q���  �@�h���h�  �PQ�҃������   �N)^�I[��_�V�   ^]� �V��+Ë^�D�����W�@��;ʋ]�E}-�F+�+�����R��R��R�I��R�x� �E��;F}L���Q���  �@�h���h�  �PQ�҃����u	[_3�^]� �N�I�ȋE�F�V)^[_�   ^]� ��U��EV���
�   ^]� W�}��|/�N;�}(�> t#�~ u%���H��0  h��h�  �҃�_3�^]� ��;�|���;���_�   ^]� S�;�|�ً�+���;��]��   ^��~�F��    QP��R�i� ���N��~;ύ��V��   ������V+���R��)F+ȉN�N�Q�+�Q�&� �F���Q���  h���h�  �PQ�҃������   �N)^[��_�V�   ^]� �V��+ÍD���~��C�^�A�;�}!�U�F+�+���Q׍�Q��R蠀 ��;^}C���H���  h��h�  ��    RP�у����u	[_3�^]� �V���F�^�])^[_�   ^]� ���U����P�B<V���Ћ��Q�M�RLj�j�QP���ҋ�^]� �������������U���VW�}���}
_3�^��]� S�]����  �F;ǋ��ύ�N�U��u(���H��0  h��hA  �҃�[_3�^��]� ��;���  )^�F�Y  @���j j�и   +�����؋F�ʙÉ]����SP�E��Â �ȉU��;�u��E�;�u�;�|�;M�r��]�Ù9U�E�|�;��{����F�U��NF�@����N��h����u���Q���  hW  P�у�����RhX  PQ��  �у��ȉ�������F�@�F�щN��~N+Ǎ@���P��+E�Í@��P��@��P�y~ +]��F����Q�[��QP�\~ ���}  �@�ҋ�+E��R�@���[R��Q�2~ ���V  ��~�N����R�@�Q��Q�
~ ���F�@��ЉN�   �F�D����@����؋F�ʙ;ʉM���   ;���   j jQS�-� �ȉU��;������E�;�� ���;E������;�������E�9U�E������;�������h����u%���Q���  �[���h|  P�у��$���J�[��h}  �RP��  �Ѓ��ȉ���s����F�@�щF�^�F;�}*�N+Ǎ@���R����E�R�@��P��| ���]�} tG�N;�}"��+��@���R�I�N��j R�{ ���V�[���P���j P�{ ���} tO�N��;�}!�F�I�Ћ�+х�t��P�P����u�V��ʅ�~�˅�t��P�P����u��؋E�F[_�   ^��]� ��������������U���VW�}���}
_3�^��]� S�]���  �F;ǋ��ύ�N�U���u(���H��0  h��hA  �҃�[_3�^��]� ��;��h  )^�F�.  @���j j�и   +�������F�ʙ��߉}���WS��~ �ȉU�;�u��E�;�u�;�|�;�r��]�Ù9U�|�;�r��M�F�V��Fы���Vh����u���Q���  hW  P�у�����RhX  PQ��  �у�����!����V�}�N���F��~>+�ɋ�+U��QӍ��Q��P�z �F+]��    Q��RP�z ���V  �ɋ�+U�Q��Q��R�mz ���7  ��~�V��    Q�R��R�Jz ���F����V�	  �F�D����@����؋F���;���   ;���   j jWS�s} �ȉU�;��A����E�;��6���;��.���;��$����E�9U�����;������h����u#���Q���  ��    h|  P�у��"���Jh}  ��    RP��  �Ѓ����������N���V�^�F9E}"�M�V+���P��P�Eȍ�Q�4y ���}�} t=�F;�}�N��+���R��j R�
x ���E�V��    Q��j P��w ���M��N[_�   ^��]� �������U����H�QV�uV�ҡ��H�U�AVR�Ћ��Q�B<�����Ћ��Q�M�RLj�j�QP���ҋ�^]���������U��Q�E;�u	�   ]� }+�RP�?���]� jj+�PR�.���]� ����������U��V��W�~��}_3�^]� jjjW�������t�F�M��_�   ^]� �������x��J| �����U��V���x��4| �Et	V�a ����^]� ���������U��M�UV�uW��r�;u��������s��tE��9+�u1��v6�B�y+�u ��v%�B�y+�u��v�B�I+���_��^]�_3�^]�����������U��QV��j �M���i �F���s@�F�M���i ^��]�������U��QVW��j �M��i �G��v	���sH�G�w����֍M�#��i _��^��]�����������������U��QW�9��t=j �M��Ci �G��v	���sH�GV�w����֍M�#��Gi ��t
��j����^_��]����U���EV�����t	V�8` ����^]� �������������̰�������������̸   �����������U��A$V�0W�}j �M�7�h �F���s@�F�M�h ��_^]� �����������U��MV3��r� ��t�����   ���ȋB(�Ѕ�u��^]� ��������������U���SVW���� �O ���EP�h P���Z� �M���  ���Q@�J$�E�PV�ы��B�P4��jh�  �M��ҡ��P�B4jh�  �M��Ћ��E�Q�R8Ph�  �M��ҡ��P�B4jh�  �M��Ћ��Q@�J(j�E�PV�ы]����3��x� ��t�d$ �����   ���ȋB(�Ѕ�u�WV����� �����   �Bj j���ЍM��/�  ���Q�J�EP�у�_^[��]� �U���4���UV��HT�Aj R�u��Ѓ��E��u^��]� S�M�Q���4� ���   +��   �]�ƨ   ���Q���������;�r��{ ���Q�F�RHW��i��   �L8 Qh�  �M��ҋN+N���Q���������;�r�{ �N��9�    _tSS���V  ���R��P�B8h�  �M��ЋM���Q�M���  ���B�P<�M�Qh�  �M��ҍM���  �M�E�P�� �M����  [�   ^��]� ������������U���L��SVW���H�A�U�R�}��Ћ��Q�Jj j��E�h��P�ы��   +��   �]�Ǩ   ���Q���������;�r�z ���Q�Rx��i��   G�M�Q���   �ҋ���H�A�ލU��R���Ѓ�����  ���QT�u�Bj	V��3Ƀ��E;�u_^3�[��]� Q�M�M�M�Qh�  �M��� P��肳 �M�躝 �����   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   �Ϋ P���V� �M��n� �����   �
�E�P�у��u�U�R���� S���T  ���Q��PP�BHh�  �M��Ћ��E�   �E�   �Q���   �E�PhT  �M��ҡ����   ��U�R�Ѓ�S���NT  ���    tUS���=T  ���Q�   P�B8h�  �M��ЋM���Q�M��R�  ���B�P<�M�Qh�  �M��ҍM���  �E�P���� �M��}�  �����   �
�E�P�у�_^�   [��]� ��������U���L��SVW���H�A�U�R�}��Ћ��Q�Jj j��E�h��P�ы��   +��   �]�Ǩ   ���Q���������;�r�;x ���Q�Rx��i��   G�M�Q���   �ҋ���H�A�ލU��R���Ѓ����T  ���QT�u�BjV��3Ƀ��E;�u_^3�[��]� Q�M�M�M�Qh�  �M�蚩 P���� �M��:� �����   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   �N� P���ְ �M��� �����   �
�E�P�у��u�U�R���9� S���1R  ���    tUS��� R  ���Q�   P�B8h�  �M��ЋM���Q�M��5�  ���B�P<�M�Qh�  �M��ҍM���  �E�P����� �M��`�  �����   �
�E�P�у�_^�   [��]� �����������U���L��SVW���H�A�U�R�}��Ћ��Q�Jj j��E�h��P�ы��   +��   �]�Ǩ   ���Q���������;�r�v ���Q�Rx��i��   G�M�Q���   �ҋ���H�A�ލU��R���Ѓ�����  ���QT�u�BjV��3Ƀ��E;�u_^3�[��]� Q�M�M�M�Qh�  �M��z� P���� �M��� �����   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   �.� P��趮 �M��Θ �����   �
�E�P�у��M�U�R�� S���P  ـ�   �5Жj �E�Ph  �M��E�   �]�E�]��Ħ P���L� �M��d� �����   �
�E�P�у�S���O  ���    tUS���O  ���R�   P�B8h�  �M��ЋM���Q�M���  ���B�P<�M�Qh�  �M��ҍM���  �M�E�P�{� �M����  �����   �
�E�P�у�_^�   [��]� ��������������U���L��SVW���H�A�U�R�}��Ћ��Q�Jj j��E�h��P�ы��   +��   �]�Ǩ   ���Q���������;�r�s ���Q�Rx��i��   G�M�Q���   �ҋ���H�A�ލU��R���Ѓ�����  ���QT�u�BjV��3Ƀ��E;�u_^3�[��]� Q�M�M�M�Qh�  �M���� P���b� �M�蚖 �����   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   认 P���6� �M��N� �����   �
�E�P�у�j �U�Rh�  �M��E�   �E�   �f� P���� �M��� �����   ��U�R�Ћu���M�Q���R� S���JM  ���    tUS���9M  ���R�   P�B8h�  �M��ЋM���Q�M��N�  ���B�P<�M�Qh�  �M��ҍM���  �E�P���� �M��y�  �����   �
�E�P�у�_^�   [��]� ����U���  �\�3ŉE�SVW���3n ��ݕ������`���ݕ�����������P�Pݝ����������Q��0���ݕ����R�荅����ݕ����3�ݝ0���P��P�����l���ݕ����ݕ8���ݕ@���ݕ����ݕ����ݝ������z�����Q�J��L���P�ы��B�PVj���L���hėQ�ҍ�L���P�N} ���Q�J��L���P�ы��   +��   �����������������d�����  ��h������   +��   ���������������9�d���r�Pp ���   �h����{ �   �}��t{���B�P������Q�ҡ��H�Ij j��U�R������P�ы�`�����������R�7[ ��\������H�A������R�Ѓ���\��� t��\���Q�5� ���U�E�RP�� ������t�������  ���   +��   ���������������9�d���r�mo ���B���   �P�h�����X���Q�ҡ��H�Aj j���X���WR�Ћ����   �R|����X���P���ҡ��H�A��X���R�Ћ��Q�J�� ���P�ы��B�Pj j��� ���h��Q�ҡ��H�U�I(R��8���P�ы����B�P��h���Q�ҡ��H�A��h���RW�Ћ��Q�J��8���P�ы��B�P�����Q�ҡ��H�I�����R�� ���P�ы��B�P<��<������ҋ��Q�RLj�j���h���QP������ҍ����P�|y ���Q�J�����P�ы��B�P��h���Q�ҡ��H�A�� ���R�Ћ��Q�J�����P�ы��B�Pj j������h��Q�ҡ��H�U�I(R������P�ы����B�P������Q�ҡ��H�A������RW�Ћ��Q�J������P�ы��B�P�����Q�ҡ��H�I��@�����R�����P�ы��B�P<��������ҋ��Q�RLj�j�������QP������ҍ����P�<x ���Q�J�����P�ы��B�P������Q�ҡ��H�A�����R�Ћ��QH���   j h�  V�Ћ��QHj �E����   h�  V�Ѓ�(�}� ǅ|���    ~g3ɍd$ �U�t��l���+���p����t+���x����t�+׉��x���+��p�P��p����P��|���B�� ��;U艕|���|���t���3�9}���   ��l���݅����݅�����M�݅�����R݅������ҋ��   ݅h�����G��܅P�����݅�����H���@����݅p����܅X���݅�����H���@����݅x����܅`������H���@�������Y��Y��Y�;}�|��������؃; �P  �}� �F  ��E�ݕ����Pݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ ���ݝ����`� ��3҃���x���;��  9U艕p�����   ��|����
�d$ ��|����M�t
���   �4v�4�V�t
�4v�4�V�t
�L
�4v�I�4���VR�������:t����   ������󥋍x���萰 ���QD��p����R0������QVP�҃�|��� F��;u艵p����i�����x�����t���j W���#� �����   �Bj j����j h�  ��诸 ����   ���Q�J��x���P�ы��B�Pj j���x���h��Q�ҡ����   �Bx�����Ћ��Q�J����,���P�ы��B�@��,���Q��x���R�Ћ��Q�B<����,����Ћ��Qj�j�WP�BL��,����Ѝ�,���Q�ot ���B�P��,���Q�ҡ��H�A��x���R�Ѓ��{ �>  ���Q�J��<���P�ы��B�Pj j���<���h��Q�ҋ��   +��   ���Q�鋋�   +��   ������������QuZ���������u�Dh ���   ����<���P���U��Q�B��W�Ћ��Q�E��JWP�у�V���k����c  ����������N  ���   +��   ���Q���������u��g ���   ����<���P���U��Q�B��W�Ћ��Q�E��JWP�у�V����������   +��   ���Q���������   �;���  ǅ|����   h)  ��� ���Q������x������~  �J������P�ы��B�Pj j�������ht�Q�ҡ��H�A(������WR�Ћ��Q�J�E���H���P�ы��B�U��@��H���QR�Ћ��Q�J������P�ы��B�P��L���Q�ҡ��H�I��L���R������P�ы��B�P<��8��L����ҋ��Q�RLj�j���H���QP��L����ҡ��H�I��<���R��L���P�ы��B�P��L���Q�ҡ��H�A��H���R�Ћ��Q�J������P�ы����   �P|����<���Q���ҋ�踤 3�9u�E�~�E�9<�u	�M�V轮 F;u�|鋍t���3��:� ��t��    �����   ���ȋB(�Ѕ�u狍t���V��x���V褳 �����   �Bj j���Ћ��   +��   ���Q���������;�r�e �����   �|�����<���R�Q���ĉE�P�B�Ћ��E��Q�JPV�ы�t�����R���9������   +��   ��|����   ���Q��������G�;��R�����t������Q�J��<���P�у���`���j j j V����L �����   �Pj j����3��������������� �������������������Ph�   �������������Cq ������   �M��l����������ą ���   +��   ��d�����h���x��������������F�d���;��D����   _^[�M�3��Z ��]ËJ��<���P�у�3�_^[�M�3��jZ ��]Í������F� �M�_^3�3�[�LZ ��]����U���SV�񋎸   +��   ���Q��������3��W�'  �]����   +��   ���Q���������;�r�c ���   E��N P�%N ����ughG  �� ��������   ���   +��   ���Q���������;�r�b �����   ���   E��R|P���ҋN j j W�J WS������WS���V����~ W��Su�����������WS���W���jj���̟ �����   �Bj j���Ћ��   +��   �E��   ���Q��������C�;������_^�   [��]Ë��B�P�M�Q�ҡ��H�Aj j��U�hؗR�ЍM�Q�Hm ���B�P�M�Q�҃�_^3�[��]�����������V�񋆈   WP��C ���   Q�C ���   �����4u  �R�\C ���   3���;�t	P�GC �����   P���   ���   ���   �&C ���N\���  �N@��  �N$��  ���Q�B��V�Ѓ�_^����U�����S�ًH�AV�SWR�Ѓ��K$蹵  �K@豵  �K\詵  j���   �@ 3Ƀ�;�t�0�3�j��N�N�N���   �@ 3Ƀ�;�t�8�3���O�O�O�Kx�K|���   ǃ�   �����F�E�9Fv�\` ��M��N�M�;Nv�G` �M��U��R�U�RQP�E�P���Ff  �w9wv� ` ��M��O�M�;Ov�` �M��U��VRQP�E�P����r  _^��[��]�����U����  �\�3ŉE�SVW��j������+�  ��,����N\P�������6�  ���Q�Bdj��,����Ћ��Q�����   h �Gh  W�Ћ��Q��j�؋BhWS��,�����j@jS�����褈  ��u+������I�������������y( u��j P�w  ��X��� �a  ���B�P������Q�ҡ��H�Aj j�������h��R�Ћ��Q�J��p���P�ы��B�Pj j���p���h�Q�҃�(������P��L���Q��������  P��p���R��<���P������P��`���Q����P��i ���B�P��`���Q�ҡ��H�A��<���R�Ћ��Q�J��L���P�ы��B�P��p���Q�ҡ��H�A������R�Ћ��Q�J��,���P�у�(��\����C�  ��\���Rǅ\������{L ��3�_^[�M�3��T ��]á��H�A��p���R�Ћ��Q�Jj j���p���h�P�ы��B�P������Q�ҡ��H�Aj j�������h�R�Ѓ�(��p���Q��������`���R跳  P������P��<���Q�C�����P��L���R�3���P�}h ���H�A��L���R�Ћ��Q�J��<���P�ы��B�P��`���Q�ҡ��H�A������R�Ћ��Q�J��p���P�у�$������B���������+  �8�����������
��$    �I ������j
������w  ��Ph�   ������Q�������  j������Rh��l �����	  ���   ���   ��������G���   ��7  �GP���H�  ������Q������hؙR�1l ���H�A������R�Ћ��Q�Rj j�������P������Q�ҋK+K���Q��������� ;�r�[ �C��������Q�RP������Q�ҡ��H�A������R�ЋK+K���Q��������ʃ�;�r�*[ �S������Ǆ�       �  j������Qhԙ�zk ����uJ���   +��   ���Q���������;�r��Z ���   �TR������h̙P�k ���A  j������Qhș�k ����uJ���   +��   ���Q���������;�r�mZ ���   �TR������h��P�j ����  j������Qh���j ����uJ���   +��   ���Q���������;�r�	Z ���   �TR������h��P�Gj ���y  j������Qh���Nj ����uC���   W����4  ��0PW���4  ��(PW���4  �� P������h��R��i ���  j������Ph����i ����uC���   W���i4  ��HPW���]4  ��@PW���Q4  ��8P������h��Q�i ���  j������Rh���i ����uC���   W���4  ��`PW��� 4  ��XPW����3  ��PP������hp�P�0i ���b  j������Qhl��7i ����uC���   W���3  ��xPW���3  ��pPW���3  ��hP������h\�R��h ���  j������PhT���h ����uV������Q������hH�R�h ��j ������P��`����O����`���Q���   W���3  �ȃ��d����`����qj������Ph@��jh ����u{������Q������h4�R�)h ��j ������P��p����AO����p���Q���   W���2  �ȁ��   �c����p������B�PQ�҃�W���2  ǀ�      ������@����������������Sk  ��u+������I�������������y( u��j P�o  j�������w�  �������^@R��膭  ���P�Bdj�������Ћ��Q�����   h �Ghe  W�Ћ��Q��jW��\���P�Bh�������Ћ�\���j@jQ��������  ��u+�������J���������������y( u��j P��n  ������ ���H�A��p���R��  �Ћ��Q�Jj j���p���h��P�ы��B�P������Q�ҡ��H�Aj j�������h�R�Ѓ�(��p���Q��`���R���c�  P������P��<���Q�������P��L���R�����P�)a ���H�A��L���R�Ћ��Q�J��<���P�ы��B�P��`���Q�ҡ��H�A������R�Ћ��Q�J��p���P�ы��B�P������Q�҃�(�������{  ���������P��������C ���Q�J��,���P�у���\����U{  ��\���R��\����C ��3�_^[�M�3��K ��]��Ћ��Q�Jj j���p���h�P�ы��B�P������Q�ҡ��H�Aj j�������h�R�Ѓ�(��p���Q��`���R����  P������P��<���Q�o�����P��L���R�_���P�_ ���H�A��L���R�Ћ��Q�J��<���P�ы��B�P��`���Q�ҡ��H�A������R�Ћ��Q�J��p���P�ы������B3���$�������������f  j
�������bn  ��Ph�   ������Q�������G�  ���   +��   ���Q��������3����   ���������Q�J������P�ы��B�@j j�������Q������R�Ћ��   +��   ���Q��������ʃ�;�r��R ���B���   ������@x������R�Ћ��Q�J���ߍ������PG�у���u2���   +��   �������   ���Q��������C�;��.����������������j������Qh$���b �����  ���   +��   ���Q���������;�r�/R ���   ��i��   ���   R������h�P�bb �������I��j
�������l  ��Rh�   ������P������蜃  ���Q�J��p���P�ы��B�@j j�������Q��p���R�Ћ��   +��   ���Q��������ʃ�;�r�uQ �����   �B���   R�P��p���Q�ҍ�p�����   j	������Qh��a ������   �������Jj
��������k  ��Ph�   ������Q���������  ���B�P��`���Q�ҡ��H�Ij j�������R��`���P�ы��   +��   ���Q���������;�r�P ���Q���   �R��i��   ���   P��`���Q�ҍ�`������H�AR�Ѓ��������A�����������3�������9�����t ����V  ��u3�������R�\_ ����t3���������������������������������������������������������������ƅ���� ƅ���� ������������������������������������������������������������������;�u)�������I��������������9y(u��WP��g  ��\���V�_ ������5  ���B�P��p���Q�ҡ��H�AWj���p���h��R�Ћ��Q�J������P�ы��B�PWj�������h�Q�ҡ��H�A��`���R�Ћ��Q�JWj���`���VP�у�<��p���R��`���P������Q��<���R������P��L���P����P��Y ���Q�J��L���P�ы��B�P��<���Q�ҡ��H�A��`���R�Ћ��Q�J������P�ы��B�P��p���Q�҃�$���H�A������R�Ѓ��������Kt  ���������Q�������< ���B�P��,���Q�҃���\����t  ��\���P��\����M< �M���_^3͸   [�_D ��]�������V�������������   ^�����������U���SVWj�0- �]3���;�t��3�jV�M��EQ�M�s�s�s�E�N8  �������   �U�U�M��+�PVQ�M��E�   �E�    �E� �IM  �U�R���N�  �}�r�E�P�. ��j�wV�MQ�M��7  �����u��UPVR�M��E�   �E�    �E� ��L  �E�P�����  �}�r�M�Q�Y. ��_^��[��]� �����������U����  �\�3ŉE�SV�uW��j������|  j@jV������xu  3���u)������H������������9y(u��WP�d  9�X����m  ���Q�J������P�ы��B�PWj�������h��Q�ҡ��H�A������R�Ћ��Q�JWj�������h�P�ы��B�P������Q�ҡ��H�AWj�������VR�Ѓ�<������Q������R������P������Q�Y�����P������R�I���P�V ���H�A������R�Ћ��Q�J������P�ы��B�P������Q�ҡ��H�A������R�Ћ��Q�J������P�у�$��\����q  ��\���Rǅ\������F9 ��3�_^[�M�3��[A ��]� ���H�A������R�Ћ��Q�JWj�������h��P�э�����R��V ���H�A������R�Ћ�����A�����������  �I j
�������d  ��Rjc������P������{  j������QhT��JZ ����uK�C|���   +��   ���   ���������������;�r�I ���   ����+��D�h�D�h�	  j������Ph����Y ����uN���   ���   +��   ���   ���������������;�r�.I ���   ����+��D�l�D�l�  j������Qh���}Y �����  ���   ���   jx�����@WR��������? ��l���   �����󥋍�������   Q����o  ���   +��   ���   ���������������;�r�H ���   ����+�3��|�d���   +��   ���   ���������������;�r�?H ���   ����+Ή|�h���   +��   ���   ���������������;�r� H ���   ����+Ή|�l3��u  j������Ph���QX �����W  �Cx�������   �������������������P�@��u�+�P������Q��������H  jj������R�������x  ������r������P�I) ��j�?' ��;�t��������������������������R�� �ĉ������������������8�p�x�� �@ ��������P�w�  ������Q軃  ������+�������$I�����������t���H����   t#��t~3���   Q���   �s!  ��d���0����   R���   �W!  ��d� ��������r  �������B  ������@������U���������ZZ  ��u)������I������������9y(u��WP�^  �{|3ɋǺ   �������Q��& ��������   h�" WjV�'>���   ���Q�J������P�ы��B�PWj�������ht�Q�ҍ�����P�$Q ���Q�J������P�у���������q  �������68  ���������R�������4 ����\�����k  ��\���P��\�����3 ��3�_^[�M�3��< ��]� 3����   3ɋǺ   �������   ���Q��% ������th�" WjV�*=���3����   ���H�A������R�Ћ��Q�Jj j�������hh�P�ы��   R������P��P��P������Q������R����P�P ���H�A������R�Ћ��Q�J������P�ы��B�P������Q�ҋ��   +��   ����������������83���r  3����   +��   ���������������;�r��C ���   ǋ@d3�@�    �������Q�$ ���   +��   ���������������������;�r�C ���   �������Tp���   +��   ���������������;�r�kC ���   ǋ@d3�@�   �������Q�2$ ���   +��   ���������������������;�r�C ���   �������T9t���H�A������R�Ћ��Q�Jj j�������h\�P�ы��   +��   ���������������;�r�B ���   �L8d�Q������R��N�����������H�A������R�Ћ��Q�R������P������Q�ҡ��P�B<���������Ћ��Q�������RLj�j�QP�������ҍ�����P�M ���Q�J������P�ы��B�P������Q�ҡ��H�A������R�Ћ��   +��   ��������������Fʃ���x;��������\����h  ��\���Rǅ\������D0 �M���_^3͸   [�V8 ��]� �����������U���  �\�3ŉE�S�]VWj���������(! 3���;�t��������������������j��������������������  ��;�t��������������������j�������������������������4q  j@jS�������j  ��u)�������H��������������9q(u��VP�'Y  9�������  ���Q�J������P�ы��B�PVj�������h��Q�ҡ��H�A������R�Ћ��Q�JVj�������h�P�ы��B�P������Q�ҡ��H�AVj�������SR�Ѓ�<������Q������R������P��L���Q�������P��4���R����P�1K ���H�A��4���R�Ћ��Q�J��L���P�ы��B�P������Q�ҡ��H�A������R�Ћ��Q�J������P�у�$�������e  ������Rǅ��������- ���������xk  �������mk  3�_^[�M�3���5 ��]� ���H�A������R�Ћ��Q�JVj�������h�P�ы��B�P������Q�ҡ��H�AVj�������h�R�Ћ��Q�J������P�ы��B�PVj�������SQ�҃�<������P������Q������R��4���P�t�����P��L���Q�d���P�I ���B�P��L���Q�ҡ��H�A��4���R�Ћ��Q�J������P�ы��B�P������Q�ҡ��H�A������R�Ћ��Q�J��t���P������ǅ���������������������ы��B�P������Qǅ���������ҡ��H�AVj�������h��R�Ѝ�����Q��I ���B�P��������@Q�ҋ������@������������  �	��$    ��j
��������W  ��Qh�   ������R�������n  j������Ph���WM ����uz������Q������h�R�M ��S��\���趑  ��\����w\P��蕕  ��\����Z�  ����  ������Q��\���聑  ��\���R���C�  ��\����(�  �  j������Ph����L �����7  ���Q�J������P�ы�������������������;�v�	< ��������������������;�v��; ������������RVSP������Q�������j  ������ǅt���   ǅp���    ƅ`��� �P�@��u�+�P������R��\�����<  jj��\���P��x����l  �   9�t���r��`���Q�D ��������R�� ���     �@   �@    �� �@ ��x�����P�u  ������Q��w  ������������+θ�$I�����������H��w��: ������9^4r�v ��� ���Q�J������P�ы��B�Pj j�������VQ�ҡ��H�I������R������P�ы��B�P������Q�ҋ��   +��   ���   ���Q���������� 3��tr�������N+N���Q���������;�r�': ���B�N������@x������R�Ѕ���  �N+N�������   ���Q��������C�;�r��N+N���Q�������   ���̍\�~  S���b  �N+N���Q���������\
��N+N���Q���������;�r�t9 ��i��   ^�Q�J������SP�ыN+N���Q���������L���������x����BǄx�����E��E��t�M��R�� ���E��     �M��    �U��    �E��     �M��    �U��    �E��e���E�    �E�ܖ��������tV���tAj �������=# �C��v	���sH�C�s����֍�����#��?# ��t
��j���ҋ�����P�E ���M��^' ��x����Q�E�Ǆx�����P�EȌ���& ���Q�J������P�у��  �����������j������Rh���nH ����u9������@P���   �������������  P������h�P�H ���`  j������QhT��H ����u:�������@���   �ЍHQ�PRP������hԚP��G ���������  j������Qh����G ����up���������   �4v�����HQP������hȚR�pG ���   ƍHQ�PRP������h��P�NG �苏�   �d�t��$��������  j������Rh���=G �����d  ���������t������P���   �b  �Ht���������������f  ������P��\�����C  jj��\���Q��x����g  ��\����2  ������R�� �ĉ0�@   �p�� �@ ��x�����P�p  ��|���Q��r  ��H�������!f  ������+�������$I�����������T����������  ���v  �#y  ��D�����������\  ��,����\  �   9������  ��    j/S��������  P��`���Q���#���P��������j  ��`����a  j �������  �xr�@���P�~F ����������NR��D�����������a  h��j�������[  P��1  ����t=j�������A  �xr�@���P� F H��������������P��,����a  ���   �v�D��ʋ���������\$�@�\$� �B�$��C;���������������������R���������$P�҃����� ������ǅ����    �w  ����������+������x�����T���ǅ����    3۹   +˃�u3ɋ�����+�P���ы������4�����������;�r��3 ���   +��   ��P����4����������������9�����r�3 ���������   �ˋ�x����Dp�����T�����+�P�������vz��<���+�8����������0��;�r�a3 ���   +��   ��8����4����������������9�����r�,3 ���������   �ˋ�x����Dp��L���T���C�������������������������A������;����������������R��r  ��8���3���;�t	P� ����,���P��8�����<�����@����~ ��P�����;�t	P�k ����D���Q��P�����T�����X����J ����  ǅ����   ���  �����������I ������j/R�������l  P��`���P������P�������g  ��`����V^  j �������9  �xr�@���P�C ��������Q���   �X��  �Pph��j�������\2���  P�.  ����t@j��������  �xr�@���P�B �X���������P���   �.  �Hp�\1������@��������;�����������������   j �������q  �xr�@���P�PB ��������������H���   R�ˉ��������  �@p������h���L0j�������  P�-  ����tFj��������  �xr�@���P��A ��������HR�ˉ������Q  �@p�������L0�������M��&#  �U�R�EȌ�� ��������3��������@�������$���3�������9�����t ����6  ��u3�������Q�V? ����t3���������������������������������������������������������������ƅ���� ƅ���� ������������������������������������������������������������������;�u)�������H��������������9y(u��WP��G  ���Q�J��t���P�ы������BǄ�������������� ǅ�������   9�����t�������5  ������Q�,> ����������������������������������������������������������������ƅ���� ƅ���� ������������������������������������������������������������������������3�ǅ����ܖ��;�tQ�8;�tBV�������� �G;�v	���sH�G�w����֍�����#��� ��t
��j����3�S�� ���������� �������H������Ǆ������Rǅ�������l ��������;�t*��|���Q������������RQP�E  ������R�j ��������P�������������������I ��������;�t*��|���Q������������RQP��D  ������R� ��������P�������������������� �M���_^3͸   [��# ��]� ���������U����  �\�3ŉE��ESV��F ���Q���   W�}j j	���Љ���Q���   j j���ЉF���Q���   j j���ЉF���Q���   j j
���ЉF���Q�J������P�у�������Rj������P����#�����Q�R�NQP�ҡ��H�A������R�Ћ��Q�J������P�ы��B�P������Q�҃�������Pj������Q���#��P��������  �������^$R���a�  �������f�  ���H�A������R�Ћ��Q�J������P�у�h���������j�  ������R���,�  ��������  ���H�A������R�Ѓ�������Qj������R����"��P�������W�  �������~@P��趃  ������軀  ���Q�J������P�ы��B�P������Q�҃�h��������  ������P��考  �������e�  j�������Z  ������Q���
�  ���R�Rhj h�   ������Q���ҡ��H�A������R�Ѓ�j@j������Q������S  ��u+������J�������������y( u��j P�B  ��h��� ���H�A�>  ������R�Ћ��Q�Jj j�������h��P�ы��B�P������Q�ҡ��H�Aj j�������h�R�Ѓ�(������Q������R����  P������P������Q蓨����P������R胨��P��4 ���H�A������R�Ћ��Q�J������P�ы��B�P������Q�ҡ��H�A������R�Ћ��Q�J������P�у�$��l����HO  ǅl�������l���R� ��_^3�[�M�3�� ��]� ������R�Ћ��Q�Jj j�������h�P�ы��B�P������Q�ҡ��H�Aj j�������h�R�Ѓ�(������Q������R����~  P������P������Q�U�����P������R�E���P�3 ���H�A������R�Ћ��Q�J������P�ы��B�P������Q�ҡ��H�A������R�Ћ��Q�J������P�ы�����J��$j
������^B  ��Ph�   ������Q������CY  ������x;  ��u+������J�������������y( u��j P��?  ������P��6 ������>  ���Q�J������P�ы��B�Pj j�������h��Q�ҡ��H�A������R�Ћ��Q�Jj j�������h�P�ы��B�P������Q�ҡ��H�Ij j�������R������P�у�<������R������P������Q������R蔥����P������P脥��P��1 ���Q�J������P�ы��B�P������Q�ҡ��H�A������R�Ћ��Q�J������P�ы��B�P������Q�҃�$�>2 ������P������������Q���b����~ t-���   +��   ���Q���������t���������/�����������1 j h  �2 ����l�����K  ��l���Qǅl������ �M���_^3͸   [�# ��]� ��������U��V��N+N��������������W�}�;�r�% �V����+�_��^]� �U��V��N+N���Q��������W�}�;�r��$ ��i��   F_^]� �����U��V��N+N��$I����������W�}�;�r�$ �V��    +�_��^]� ���������������U��V��襥���Et	V�9 ����^]� ��������������̡�V��H�QV�����V ���   �V(R�V0�V8�V@�VH�VP�VX�V`�Vh�Vp�^x���H�A�Ћ��Q�J���   P�ы��B�P���   Q�ҡ��H�A���   R�Ѓ���^á�V��H�A���   R�Ћ��Q�J���   P�ы��B�P���   Q�ҡ��H�A���   R�Ћ��Q�BV�Ѓ�^��������U��V��V����� ���Et	V�� ����^]� �����U��A�U��Q �E��U+ЋA0�]� ��������������̋A �8 t�I0��3�����������������U��A�U��Q$�E��U+ЋA4�]� ���������������V���F@t�F�Q�\ ���V�    �F �     �N0�    �V�    �F$�     �N4�    �f@��F<    ^������̍Q�Q �Q�Q$�A�A�Q(�Q0�A�A�Q,�Q4�     �A$�     �Q4�    �A�     �Q �    �A0�     ���������U���SV��H�QWV�ҡ��H�}�QVW���G�^���   �GS�^�G�F�O �N �W$�V$�G(�F(�O,�N,�W0�V0�G4�F4�O8�N8�W<�V<�G@�F@�OD�ND�WH�VH�GL�FL�OP�NP�WT�VT�GX�FX�O\�N\�W`�V`�Gd�Fd�Oh�Nh�Wl�Vl�Gp�Fp�Ot�Nt�Wx�Vx�G|�F|���Q�B�Ћ��QS���   P�J�ы��B�H���   S�ы��B�P���   SQ��ه�   ٞ�   ���H�Q���   S�ҡ��H�A���   SR�Ћ��Q�B���   S�Ћ��Q�J���   SP�ы��   ��<_���   ��^[]� ��������U��VW�����u�  ���t��3ҋE����+��G����;Bw��t�	�3�;As�� w��_^]� ���������U��VW�����u� ���t��3ҋE�4�    +��G���;Bw��t�	�3�;As�{ w��_^]� ���������U��M����w3ɋ���+����R�.�  ����]Ã��3����xsڍEP�M��E    �� h���M�Q�E�x�� ���U��M����w3�i��   Q���  ����]Ã��3���=�   sߍEP�M��E    �r h���M�Q�E�x�� ��������U��M����w3ɍ�    +���R�n�  ����]Ã��3����sڍEP�M��E    � h���M�Q�E�x��Z ���U��M����w3ɍ�    R��  ����]Ã��3����s��EP�M��E    � h���M�Q�E�x��  ���������U��EVP���� �x���^]� ����U���VW�}��H�QVW���G�^�G�^�G�F�O �N �W$�V$�G(�F(�O,�N,�W0�V0�G4�F4�O8�N8�W<�V<�G@�F@�OD�ND�WH�VH�GL�FL�OP�NP�WT�VT�GX�FX�O\�N\�W`�V`�Gd�Fd�Oh�Nh�Wl�Vl�Gp�Fp�Ot�Nt�Wx�Vx�G|�F|���Q�R���   P���   Q�ҡ��H�I���   R���   P��ه�   ٞ�   ���B�@���   Q���   R�Ћ��Q�R���   P���   Q�ҋ��   ��(���   _��^]� ���U��S�]V�u;�t#W�}V���������   ���   ;�u��_^[]ËE^[]��������U��S�]V�u;�t#W�}���   ���   V���I���;�u��_^[]ËE^[]��������U��E��V��M�Q�F����� ��V�H�N�P�V�@�F����^��]� ���������������U���E��QP�p ��]� ��������U��S�]V�u;�tW�y�WP�D �F��;�u�_��^[]� U���E��QP�|
 ��]� ��������U��S�]V�u;�tW�y�WP�P
 �F��;�u�_��^[]� U��E]� ������U��E�UV�1W��+�W�}WP�FR��_^]� �������������U��S�]VW�}��+�9us� �E�MVSPQ� ����_^[]� �����������U��E]� ������U��E�UV�1W��+�W�}W�}WP�F(R��_^]� ���������U��S�]VW�}��+�9us�- �E�MVSPQ�- ����_^[]� �����������U��V��F�����~�FP�G �}�NQ��  ���E���t	V��  ����^]� �������̃��� ����������3��������������̃���������������U��U��@R�Uj�R��]� �������̋�� ������������ ������������̋A$�8 t�I4��3����������������̋A �8 t�Q0�: ~� � Ë�B�����V���P�҃��u�^ËF0��F ��Q��^����������U��E����3ɉH�H�H]� ���U��E����3ɉH�H�H]�  ���U��A � ��t<�Q;v5�U���t:P�t�A@u"�A0� �A ����t�A ����]� 3�]� ���]� ̋Q V�2��u���^�SW�y0����;�s�_[^��A@u/�A$� ��t&;�w9q<v9A<s�A<��A<+�I ��_[^�_[���^����������������U��SV�q$�W��t9A<s�A<�]����   �A �����   �E��u�A�y<+8�u��'��u��u�A�u��+8����t�5����u����   �A� �y<+�;���   +Q0�)�Q ����   �Q$�����   �Q4�ЋA R��AR�R�[����p��te���t_�E�=����u�A�Y<+�u����u�A�u��+��	����u�u��|�A� �Y<+�;�+Q4�)�I$�
����5���E_3ɉ0^�H�H�H[]� ��U��E�UVW�y$�4���t9A<s�A<���;���   S�]$��tR�Q ���tI��|w�A� �y<+�;�d+Q0�)�Q ��tX�Q$���tO�Q4�ЋA R��AR�R�K����4��t-�?��t'��|#�A� �Q<+�;��Q4+��)�I$������[�E3�_�0�H�H�H^]�  ��������������U��V�q���Q�F�D���P� ���; ���Et	V�^�  ����^]� ����U��V��W�~8�ܖ��t��蕖��W�/�  ���N�H �Et	V��  ��_��^]� �������������U��V��W���~����~8�ܖ��t���:���W���  ���N�� �Et	V��  ��_��^]� ��U��Q�U�E�M���u	;A��   SVW�y;�st+�;�wn�   +���yr
���M�	����M��E�WQS� ������t5�U�ERPV蟔������t,�M�+ލ|�WR�^S�� ������u�_^���[��]� �E��x�Mr�	_��^+�[��]� �U��SV�uW��9ws�� �G+Ƌu;�s���]��;�r�Ãr�����MP�EP�W��������u;�s
_^���[]� 3�;���_^[]� �U��M����w3�Q�k�  ����]� ���3����s�EP�M��E    � h���M�Q�E�x��U �������������̋A �8 t�Q0�: ~����I ��P�� Ë�P���������V�����t(��u�� ��xr�H��H�@�9Fr�� �F^����������U��E��u&�yr�I�E�U�]� �E�U���]� �yr�I����UP�EP�Q�p	 ��]� ���������U��QS��V�K�ܖ�D j�3�  ������t@W�� ��� j �M������ �G���s@�G�M���� _�ˉs8�����^��[��]�3��ˉs8�����^��[��]�������U��S�]V�uW���    ��t)��t%�V�F��r����;�w��r� �N�;�v� �7�_��_^[]� ������������U��E�M�UV�uPQRV�} ����^]����������������U��E�M�U ��E��   ]� ����U��E�M��   ]� ������������U��E+E�M;�s��]� ����������U��S�]V�u��+θ����������������+ȋE�ȉM��;�t#+�W��I �<���x�   �;�u�E_^[]�^��[]����������������U��W�}��tV�u�   �^_]� ����U��M��t	�EP����]� ���������U��S�]V�u��+˸����������������+���ɋыM��+�;�t+�W�M��M��x�<�   ���;�u�_^[]����������������U����US�]V�uW�}2��E��M��E��E�PQRWVS�r���+���Q���������i��   ����_^+�[��]����������U��j�h��d�    PQSVW�\�3�P�E�d�    �e��E�    �]�}�u��$    ;utVW��������x�}��x�u���E������ǋM�d�    Y_^[��]�j j � ����������������V��F � ��t=�N0�	��~�F0��F � �V �� ^Å�t�N0�9 ~����F ��Q���	��P���҃��u�^ËF �8 t�N0�9 ~��^Ë�P��^������U��QV3�9uW���u�~nS�]���s�����~6�M;ȋ�}��G ��UVQRS�9 �G0)0u�)u�G ރ�0�u����P���҃��tF�C�M�u��} �[_��^��]� _��^��]� ������U��QV3�9uW���u�~mS�]���s�����~3�M;ȋ�}��VSP�G$�Q�
 �G4)0u�)u�G$ރ�0�u����P�B���Ѓ��tFC�M�u��} �[_��^��]� _��^��]� ������̋A��PV�q��D
��W���������~8�ܖ��t���\���W���  ���N�� �F��H_�D1���^�����������U���V���F@Wt �~$���t�N<;�s�F4� +��N4��E���u
_3�^��]� �V$�:S��t$�N4����;�s�	�v$�[�Q�_�^��]� �F@u=��u3���F4�N�+ߋ���� s�    ���v������+�;�s��u��u[_���^��]� �P�ND�E��������F��M���vSQ�M�QW�y����M�����u"�V�~<�:�F$�8�V4�E���F@u7�GPW�V�F$��+�V<� �V��+�+��V$ǉ��+�U��F4��F@t�V�:�F �     �V0�:��F$��F BR�+��RW���o����M��F@t	Q�P�  ���F4�N@��v$��A��E[_�^��]� ������������U��S�]V��W9^s��� �F�}+�;�s����v^�N��r�V��V�U��r�V��V+�P�E��P+�Q�R� 	 �F+ǃ��~�Fr�N_� ��^[]� �N� _��^[]� ��U��} VW�}��t'�~r!�FS���vWSjP� ��S�]�  ��[�~�F   �D> _^]� ����U��E�MPQ� 3҃������]�V��~L t#��Pj��҃��t�FLP�� ����}���^�3�^�U��A � S�]��t,�Q9s%���t�@�;�u�A0� �I �	��@���#�[]� �AL��t$���t�y< u��PQ� �����t��[]� ���[]� �V��F ���t�Ћ�V0��;�s�^Ë�PW���ҋ����u_�^Ë�PW���ҋ�_^������������U��V��NLW��tl�U�}��u	��u�G�3�WPRQ�D ����uG�~L���FH�FA�������t�G�F�F�G�~ �~$�F0�F4�~L���FD_�F<    ��^]� _3�^]� ��������������U��ES�]V���F<    �F@����   ��<tzWS�ND��������ESPSW� ���F@��F<u�N�9�V �:�N0��N@��u7��u�ǋV�:�N$���+ЋF4Ӊ�N �9 u�V�:�F �     �N0�9�N@_^[]� ����������U��V�1W�y��u�� 3��Mi��   �;xw��t�����3�;xs�� �E�x_�0^]� �����U��j�h��d�    P��SVW�\�3�P�E�d�    �e����}�E�������v���"�_���鸫�������;�s�����+�;�w�4�E�    �NQ�������؉]��E������0�e��E�E�E�@P�M������E��E�   ��Ë}�u�]�M��v �r�G��GQP�VRS�� ���M�r�GP��  ���M�G�  ��w�O��r��� �M�d�    Y_^[��]� �u�~r�NQ�r�  ���F   �F    �F j j �{ ����U����US�]V�uW�}2��E��M��E��E�PQRWVS�����+���Q���������i��   ���_^[��]��������������U��E�U;�tS�]VW����x�   ���;�u�_^[]�������U��V�uW�};�tS�]S����������   ;�u�[_^]�������U��E�M;�t�UV�2�0��;�u�^]��U��j�h��d�    PQSVW�\�3�P�E�d�    �e��E�    �]�}�u��$    ��v�EPV������O�}��x�u���E������M�d�    Y_^[��]�j j � ��U��j�h �d�    P��SVW�\�3�P�E�d�    �e��}�}��E�    �]�u��;utVW���R������   �}���   �u���E������ǋM�d�    Y_^[��]Ëu�};�t����������   ;�u�j j �v ���������������V�qP������V������ ��^�����V��~r�FP��  ��3��F   �F�F^�����������U��VW�y��wP������V����� ���Et	W���  ����_^]� ��������U��yr�AV�uQP���������^]� V�u�AQP��������^]� ���������U��V�������E3����u�   �u���t���t���E�x�Pr�@QRP��������^]� Q��RP���o�����^]� ��������U��U��V�p�d$ �@��u��M+�P�ARPj ����������^]���������������U��Q�M�U�E� �E�P�EQ�MR�UPQR�k�������]�����U��Q�M�U�E� �E�P�EQ�MR�UPQR��������]�����U��j�h �d�    P��SVW�\�3�P�E�d�    �e��u�u��E�    �]�}����v�EPV�������O�}���   �u���E������M�d�    Y_^[��]Ëu�};�t���G������   ;�u�j j �� ���̃y$r�AÍA���U��V���H��~$r�FP��  ��3��F$   �F �ΈF��� �Et	V�p�  ����^]� ������U��V���T��~$r�FP�E�  ��3��F$   �F �ΈF�� �Et	V� �  ����^]� ������U��SV3�S���� �^�   �F�^�F8�^4�^$�FT�^P�^@�Fp�EP�^lV�^\��� ����^[]� ���SV��WV�L� ���~pr�F\P��  ��3ۿ   �~p�^l�^\�~Tr�N@Q��  ���~T�^P�^@�~8r�V$R�f�  ���~8�^4�^$�~r�FP�K�  ���~�^_�^��^[�� �����U��S�]V�����+F;�w��� ����   W�~����v�� �F;�s9�NQW���L�����vZ�U�FRSP���(����~�~r:�F�8 _��^[]� ��uщ~��r�F_�  ��^[]� �F_�  ��^[]� �F�8 _��^[]� �����U��S�]VW�}��9_s�N� ��E+�;�s���M;�uj��W���'���Sj ������_��^[]� ���v��� �M�F;�s�FPW���t����M��vj�yr/�I�-��u�~��r�F_�  ��^[]� �F_�  ��^[]� ���~�^r���ËUW�Q�NQP��� ���~�~r��; _��^[]� ����������U��USVW���tF�~�F��r����;�r1��r���ȋ^�;�v��r� �MQ+�RV�������_^[]� �}���v��� �F;�s�VRW���{�����vY�N�^��r.��,��u�~��r�F_�  ��^[]� �F_�  ��^[]� �ËUWRQP��� ���~�~r��; _��^[]� �����U��Q�UV�uW�}�E� �E�P�ER��QPVW�����΃���+΍�_^��]� ����U��V3���j��F�F   P�F�EP�������^]� ��������U���D�\�3ŉE��A �8 �M�t/�Ћ�Q0��;�s �A0��A ��Q���M�3���� ��]ËAL��u����M�3���� ��]Ãy< uP� �����t����M�3��� ��]�SVWP�E�   �E�    �E� � ������  ��Pj�M��U����}��E���A  ���u؅�t!�ȃ�s�M�;�w�ȃ�s�M�U��;�v�^� �}��U�E�M����t�ȃ�s�M��;�r�8� �}��U�E�ڃ���   ����t�ȃ�s�M�;�w�ȃ�s�M��;�v��� �}��U�E�M����t��s�E��;�r��� �}ЋO<��R�E�P�E�P�E�P�E�P�E��PV�GDP�҅��   ��~k����   �}���   j�U�R�M��������s���P�E�jP�}� �u߃��M��(���_��^[�M�3��.� ��]ÍM�M؋������u������E�9E���   �U��E����   ����t!�ȃ�s�M�;�w�ȃ�s�M�]��;�v��� �U��E�M����t��s�E�U��;�r��� �E�+�Pj �M������OLQ�� ������ ����M��h���_^���[�M�3��m� ��]Íu��m����}�M�Q�M��������f���+}ԋ����~�UЋBL�M��T�NPR� ������uߍM������M�_��^3�[�� ��]����������������U��V�u��W�x�I �@��u�+�PV�P���_^]� ����������U��SVW�}���    ��t�E9Fw;Fv��� �E�]���G9^w;^v�� �]����t;�t�� �O;�t!�F�E �UR�UR�URQPS�w������F��_^[]� ��������U���,�\�3ŉE��y< �M���  �yA ��  ��Pj��҃��u2��M�3���� ��]ù   3��E� �M��E�E��E�   ��s�E�SV�@ W�E�U����  �؉]؅�t!�ȃ�s�M�;�w�ȃ�s�M�u��;�v�� �U��E�M����t�ȃ�s�M�u��;�r�� �U��E�}����   ����t$�ȃ�s�M�;�w�ȃ�s�M�]�ˋ]�;�v�C� �U��E�M����t��s�E�U��;�r�� �E܋H<��R�E�P�E��SV��DP�҃� t<��t>���M��R  ����_^2�[�M�3��� ��]Í]�]�������u��V����E��@A �U��E����   ����t!�ȃ�s�M�;�w�ȃ�s�M�}��;�v�� �U��E�M����t�ȃ�s�M�}��;�r�Z� �U��E�}�+�tv����   ����t!�ȃ�s�M�;�w�ȃ�s�M�]��;�v�� �U��E�M����t��s�E�U��;�r��� �E܋HLQWjV�m ��;�u7�U��E�M܀yA t0�������Wj�M��t���������u������u��h����M������M��_���_^�[�M�3��e� ��]ËM�3Ͱ�U� ��]�������������U��V�uW�}�Ƌυ�v�US��H����w�[��_^]� ���U��V�uW�};�t����y������   ;�u�_^]� ���������U��Q�UV�uW�}�E� �E�P�ER��QPVW�i�����i��   ���_^��]� ����U��Q�U�E� �E�P�ER�U��Q�MPQR�+�������]� ��U��V�u�~r�FP�j�  ��3��F   �F�F^]� ���U��S�]V�u;�t!W�}j�j V����������;�u��_^[]ËE^[]����������U����\�3ŉE����M;�tT�PS�XV�p�]��YW�x�X�Y�X�Y�X�Y�X�Q�U��q�q�y�Q�P�p�q�Q�P_�p^�Q[�M�3��� ��]� ���U��V���9� 3��N�H�j��A�A   P�A�EP�������^]� ����������U��V����� 3��N�H�j��A�A   P�A�EP�����`���^]� ����V���H��~$r�FP���  ��3��F$   �F �F��^�S� ��������������U��V�u3�j��NQ���F   �NP���*�����^]� ���U���   SW�}3ۉ]���tm9uiVj�}�  ������t)�Mj �E�P�   ����P��l����E���P���m����3��^��t��l�������s�����t�}�r�M�Q��  ��_�   [��]��U��V���� 3��N�T�j��A�A   P�A�EP�a����l���^]� ����V���T��~$r�FP��  ��3��F$   �F �F��^�� ��������������U��UV���W�F   �F    �F �x�@��u�+�PR�������_��^]� �����U���4�\�3ŉE�S�]�щU܃��u3�[�M�3��� ��]� �J$�9 Vt/�B4�	�0�;�s"��B$��Q��^��[�M�3���� ��]� �BL��t�z< u'P��P�� �����u�^���[�M�3��� ��]� �   3��E� �]؉M��E�E��E�   ��s�E��@ W�E�U������  �؉]ԅ�t!�ȃ�s�M�;�w�ȃ�s�M�u��;�v�_� �U��E�M����t�ȃ�s�M�u��;�r�9� �U��E�}����  ����t$�ȃ�s�M�;�w�ȃ�s�M�]�ˋ]�;�v��� �U��E�M����t��s�E�U��;�r��� �E܋H<��R�E�P�SV�E�P�E�P�E�P�E܃�DP�҅���  ���A  �U��E���"  ����t!�ȃ�s�M�;�w�ȃ�s�M�}��;�v�`� �U��E�M����t�ȃ�s�M�}��;�r�:� �U��E�}�+�tz����   ����t!�ȃ�s�M�;�w�ȃ�s�M�]��;�v��� �U��E�M����t��s�E�U��;�r��� �E܋HLQWjV�M� ��;���   �U��E�M��AA�M�9M���   �������}� �M���   j j�;���������]�]�������u��I����u�������u��<�����uu�U܋BL�M�PQ���������t �u�M������_��^[�M�3��� ��]� �M���������_��^[�M�3���� ��]� �M������E_^[�M�3���� ��]� �M������M�_^3̓��[�� ��]� �����������U���SV��F W�~@98u�}u�~< u�]K��]�~L ��   �'�����tw��u�}t�M�VLQSR�e� ����uX�NL�E�PQ�Y� ����uD�V 9:u�N�9�V �FA�Ή�V0+ȃ�A�
�E�M��U�_�H�ND^�     �P�H[��]� �E���_3�^��H�H�H[��]� �������������U����EV��~L �MW�}�E��M���   ���V�����t�FL�U�RP�$� ����uk��t�NLjWQ�� ����uT�FL�U�RP�|� ����u@�M�V �ND�N@9
u�FAPPQ���F����E�M��U��H�ND_�     �P�H^��]�  �E���_��@    �@    �@    ^��]�  �����������U��QSVW�}���    ��t�E9Fw;Fv��� �E�]���G9^w;^v�� �]����t;�t�� �G;�tB�VPRS�&����؋F���E���;�t��I ����������   ;}�u�E_�^^[��]� ��_^[��]� ����S��V�s3�;�t(W�{;�t���������   ;�u�CP��  ��3�_^�C�C�C[����������������SV��3�W��9^Lt������u3��FLP�� ����t3��Έ^H�^A�����^L����_�^<�ND^[����U��VW�}W���� 3�j��N�H��GR�A   �QP�Q�����_��^]� ����U���DSj3�ht��M��E�   �]��]������M���� j�S�E�P�M��E�H��E�   �]܈]�����h(��M�Q�E�`��� �����������U��VW�}W����� 3�j��N�H��GR�A   �QP�Q�,���_�`���^]� ��������������U���SVWj �M��5� �=� ���]�u+j �M��� �=� u��@�����M�� � �}�5��;ps"�H����u�x t�� ;ps�P�4��3�����u]��t�M����� _��^[��]ÍE�WP�C��������uh���M��f� h���M�Q��� �u��Ή5��j��V�� ���M��� _��^[��]�������U��Q�U�E� �E�P�ER�U��Q�MPQR�{�������]� ��U���   SW�}3ۉ]���tp9ulVj�=�  ������t,�M�E�P�   �S���P��l��������F    �T��3��7^��t��l�������0�����t�}�r�M�Q���  ��_�   [��]���������������U����US�]V�uW�}2��E��M��E��E�PQRWVS�B���+�$I�������������    +ȍ�_^[��]��������U��V�uW�};�t*S3ۃ~r�FP�?�  ���F   �^�^��;�u�[_^]����U��M3�;�tj��A�A   P�A�EP�{���]� �������U��j�h@�d�    P��SVW�\�3�P�E�d�    �e��}�}��E�    �]�u��;utVW���������}���u���E������ǋM�d�    Y_^[��]Ëu�};�t�]V���������;�u�j j �{� ����U��E���A�I��D#���   �} t	j j �N� ��t'hĘ�M������E�P�M������h��M�Q�"� ���M�t$h���Y����U�R�M������h��E�P��� h���5����M�Q�M�����h��U�R��� ��]� �����U��VW�}W���� 3�j��N�T��GR�A   �QP�Q�����_��^]� ����U��VW�}W���h� 3�j��N�T��GR�A   �QP�Q����_�l���^]� ��������������U��QS3�V��WSS�^$�^�^�F  �F   �^�^�^ ����j���  ����;�t6�/� ��V� j �M����n� �C���s@�C�M��� �~$_^[��]�_�^$^[��]���������������U��V��~H ��t����W�~8�ܖ��t���f��W�N�  ���N�g� �E_t	V�6�  ����^]� ������������U����A$SVW�8j �M��}��� �G���s@�G�M���� �M�Q�X�����j �M����� �G��v	���sH�G�w����֍M�#��� ��t
��j���Ћ�E�RP����_^[��]� ��U��V3�W�}��F�F�F;�u_2�^]� ��I�$	v����PW���������    +ύ��F�F_�V�^]� �����������U��j�h`�d�    P��   �\�3ŉE�SVWP�E�d�    �e��ًC��u3���K+ȸ���������������} �i  �s��p�����+K��������������º"""+ЋM;�s�L����;��,  ����"""+�;�s3���;�s��j W�������ȉ�p����u+s����������������E�    �EP�UR����+ƍ�Q���z���ǅl���   ��p���R�EP�KQ���Z���ǅl���   �U����+Ƌ�p�����R�CP�MQ���+����E������s�K+θ��������������E��t	V��  ������+ϋ�p����ȉS�M����+эЉK�C�  ��p���R�r�  ��j j �� ��+M��������������¹   �u��t����;E��   �}����+�����E�Q��p���RP���_����E�   �K��t���P+M���������������+�W�CP���*����E�����s�[��t���R+�S�EP��������N�E����+������p�����+�PPW��������C��p���QW�UR������t���P�E�VP�z������M�d�    Y_^[�M�3��D� ��]� ���������U��j�h��d�    P���   SVW�\�3�P�E�d�    �e���u�F��u3���N+ȸ��Q��������ڋ}����  �N��+V���Q��������º�G+�;�s�h����8;��g  �����G+�;�s3���;�s��j S�������ȉM�U+V���Q��������E�3҉U��U��URWi��   �P���[����E�   �E�P�MQ�VR�������E�   �E��i��   E�P�NQ�UR���|����E������N�V+Ѹ��Q������������t�VRQ�������FP���  ��i��   �E�؉^i��   ��~�F�M�d�    Y_^[��]� �]��u�}��~��i��   �QW�M��\�����~ �U�i��   �Pi��   �V�M��8���W�R�  ��j j �m� +M���Q���������;ύ������   �UR�k�����i��   �E�Q�VRP���p����E�   �N�����P+M���Q���������+�W�FP��������E�����^�v�����R+�V�EP��������p�Ei��   �M�Q�R�U�P�k���j j �� �EP�ɼ���^i��   ��+ǉESSP��������FS�MQ�UR���������P�E�WP�{����������蝺���M�d�    Y_^[��]� ���������U��j�h��d�    P��SVW�\�3�P�E�d�    �e���V��u3��
�F+����ȋ}����  �^��+�������?+�;�s�Y����8;���   �������?+�;�s�E�    �M��ȉM�;�s�U��j Q�=������E�]+^���E�    �MQW��R��������E�   �EP�MQ�VR���#  �E�   �;�]��Q�VR�EP����"  �E������F�N+������t	P��  ���U���F���N�^�M�d�    Y_^[��]� �UR轾  ��j j ��� �ˋE+���;�sv�U�
�M��    �M�QSP���e"  �E�   �F�UR��+M��+�WP�������E������EF�v�UR+�V�EP�������M�d�    Y_^[��]� �M��U��    �E��+�SSW����!  �FSW�EP�!  �MQ�E�U�RP�\������M�d�    Y_^[��]� �����U��Q�M�U�E� �E�P�EQ�MR�UPQR���������]�����U���SVWj �M��E� �=� ���]�u+j �M��)� �=� u��@�����M��0� �}�5��;ps"�H����u�x t�� ;ps�P�4��3�����u]��t�M����� _��^[��]ÍE�WP���������uh���M��v� h���M�Q��� �u��Ή5��[��V�� ���M��� _��^[��]�������U��V�uW�};�tS�]j�j S��������;�u�[_^]������U��j�hЊd�    P��SVW�\�3�P�E�d�    �e��u�u��E�    �]�}����v�EPV��� ���O�}���u���E������M�d�    Y_^[��]Ëu�};�t�]V���f�����;�u�j j ��� ������U��E�MP����]����������������U��U��t�Ay( u���URP�>���]� ���������̋A��PV�q��D
����~H W��t���z����~8�ܖ��t���Z��W�@�  ���N�Y� �F��H_�D1���^�����U��EVWP���p�������B�����Є�t�G<    _^]� �ωw<�׶��_^]� �Vj���ָ  3Ƀ�;�t�0��N�N�N��^�3���N�N�N��^������������U���   �\�3ŉE�SV�ًCW�   �u�}��{�u��+ȸ��������������;�vH9{v�d� �K+K�E�P���������������+�VWP�������_^[�M�3��
� ��]�| s]9{v�� �K���t����M�;Kv�� �M���M�V��|�����|����������t����M���|���WPQR��t���P��������M�_^3�[�� ��]�| �������������U���SV��^�F��+ȸ��Q��������W�}�;�vD9^v�p� �V+V��EP���Q���������+�WSQ��������M蘳��_^[��]�� sN9^v�*� �F��M��E;Fv�� �E��E�W�E�P�M��U�������M��P� SQRP�M�Q��������M�7���_^[��]�� ��������������U��E�UP��Q�MQR�8�����]� �U��V��~L W��   �E�M�UPQR�a� ��������   ���FH�FA �B����N8�G�F�F�G�~ �~$�F0�F4�~L���FD�F<    �9j �M�}��� �G���s@�G�M��� �UR�Y�������P�����҄�t�M�F<    �8W��_��^]� �Ή~<足���M�W��_��^]� _3�^]� ��������������U���SV��FW�~��+�������u3��#;�v�� �M���t;�t�{� �]+����U�E�MRjPQ���7����~;~v�Q� �6�u��}���u�@� 3��<�;xw��t�6����3�;~s�� �E�U��x_^�[��]� ���U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U��j�h��d�    P��0�\�3ŉE�SVWP�E�d�    �e��}�u�ủu��E�   3��E�EԉE��]�;}t$�E�PV���?���WV���������ũ��}����E������}�r�M�Q�1�  ���ƋM�d�    Y_^[�M�3��	� ��]Ëuȋ}�;�t�]�I V���x�����;�u�3�PP�� ��������V���HW�13��@u�@(��ȋB0�Ѓ��u�   ��I΅�t�Aǃy( u��j P�E���_��^�U��QV��F��t�M�Q�N�VRQP�����VR�g�  ���P�F    �F    �F    �G�  ��^��]����������������U���V��NW��u3���F+����~��+���;�s�E�����~_^��]� ;�v��� �U�RWP�E�P���4���_^��]� ������������U��VW�y��wX���.���V����p� ���Et	W蓴  ����_^]� ��������U��j�h �d�    P��SVW�\�3�P�E�d�    �e���u��H΋A����   �I,��t�R����} up��P�L2��tb�MQ����T��P�{��������M�^S���E�    ��B�L0(�ٸ���E���uj j��I��!�����ЋG�PHu+�E�������Q�2�y ue��M�d�    Y_^[��]� ��Q�L2(����럋M��@��H���x( u�����H�Hu�E������9GËu��j j �p� �A���y( u��j P�����2��M�d�    Y_^[��]� ������������U��SVW�}���    ��t�E9Fw;Fv� � �E�]���G9^w;^v��� �]����t;�t��� �O;�t5�F�E �UR�UR�URQPS������V�؋EP�NQRS�#�����(�^��_^[]� ����U��Q�UV�uW�}�E� �E�P�ER��QPVW���������    +΍�_^��]� ��U��SV�uW�}��+ϸ�$I�����������    +ȋE�ɋ�+�;�t+ƉE��E��V�0�����;�u�_^��[]�����U���SV��FW�E�9Fv��� �~�;~v�� �M��QSWP�U�R������_^[��]������������U��QS3�VW�ىE�9Et���CX����Q����C��p���3����{j �Ή~(�F,    �����~( �F0u�F��j P��������F    ��Q�����誼�������GH �GA �լ��3��GL���G<�OD_^��[��]� ���������U��QS3�VW���E�9Et���GP����Q����G��p����s����_j �Ή^(�F,    �M����~( �F0u�F��j P�������E�F    ��Q�M��PQ����������_^[��]� ����U��j�h@�d�    P��SVW�\�3�P�E�d�    �e���u�3ۉ]�^�u܋�H�D1(;�t�H�� j���G�����tY�}��~R�E�    ��B�L0(藴���E���u���&�M;�u�F��Q�L2(�a����O�}��m���]��E������E�  �~ u���Ӌ�I΅�t�Ay( u��j P������E܋�J�D(��t�H�d� �ƋM�d�    Y_^[��]� �F�M�A�M��H�L1(� ����D����M��B��H���x( u�����H�Hu�E�������KËu�]��E���j j ��� ������U��j�h`�d�    P��$SVW�\�3�P�E�d�    �e�3��}��E� �u�uЋ�H�D1(��t�H茻 j �����������   ��BƋ@$�8�}�j �M��߶ �G���s@�G�M��� �E�P�z������E܍M��\M��j�j �]��������E�    ��Q�2�A��~���r��������}؋I(豲���E��v	���uq�M��E������}��H�D1    �}� u����J΅�t�Aǃy( u��j P� ����EЋ�Q�D(��t�H蜺 �ƋM�d�    Y_^[��]��ȋU܋R�JHu�Pj��������E�O�}؋�H�L1(�E����O����M��B��H���x( u�����H�Hu�E�������MËu�-���j j ��� ��������������U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U��Q�M�U�E� �E�P�EQ�MR�UPQR�;�������]�����U��QVW�}��;��W  �G�O+ȸ�$I����������Eu���V���_��^��]� �NS�^+˸�$I�����������9MwY�GSP�GP�����MQ�N�VRQP�{����O+O��$I�������������    +ЋF[��_�N��^��]� ��u3���V+ӉU���$I���U��������9Ew+�G��    +э�SQP�M�����F�O�U��PQR�M��t�FPS�������FP�5�  ���O+O��$I�����������P��������t�N�W�GQRP���
����F[_��^��]� ������������U��j�h��d�    P��<�\�3ŉE�SVWP�E�d�    �e���u��E�E��F��u�E���N+ȸ�$I����������E̋}����  �^��+N��$I����������¹I�$	+�;�s�����ǋM�;���  ����I�$	+�;�s�E�    �M��ʉM�;�s�E̋�j Q�|������ȉMȋ]+^��$I����������ډ]�3��E��E��U�RW��    +Í�Q���W����E�   �U�R�EP�NQ��������E�   ߍ�    +ӋEȍ�Q�VR�EP��������E������^�N+˸�$I��������������t�VRS�������FP�H�  ���E̍�    +ȋEȍ��V��    +ύ��V�F�  �]��uċ}ȃ�~��    +ƍ�QW�M��E�����~(�U���    +ȍ�R��    +ƍ�Q�M�����W�è  ��j j ��� +]��$I�����������;���   �M�Q�M�������    +��ۋE�R�NQP�������E�   �N�U�R+M��$I�����������+�W�FP��������E�����^�v�M�Q+�V�UR�~������~�M��    +����M��Q�R�U�P�E���j j �� �E�P�M��p����F�Eč�    +��ۋ�+�PPW��������F�M�QW�UR�����E�P�E�SP��������M��s����M�d�    Y_^[�M�3��p� ��]� �����U��EV���F�@   �@    �@ ���t#PQ������Q���D��t�    ^]� ��^]� U���SV��^W�~��+ϸ�$I�����������u3��3;�v� � �M���t;�t��� �M+ϸ�$I������������M�U�EQjRP��������^;^v�� �6W�M��u��]��ܤ���E�M��U�_^��P[��]� �����U���SVW���G��u3���O+ȸ�$I�����������_��+O��$I�����������;�s.�U�E� �M�Q�MR�GPQjS���������__^[��]� 9_v�� �U�RSP�E�P������_^[��]� ���������������U��EW�};E,tQ���u�� �ML�EP�+����E��u�� �E��t#�MQP�������J���Dt3��E��E;E,u��}(�UL�r�EP�L�  ���}H�E(   �E$    �E r�M4Q�(�  ����_]�U��QSV�u3ۈ]��E��M��U�P�ELQ�M,RP�� �ĉj��HS�U0�A   �YR�Y�\����M�� �ĉj��HS�U�A   �YR�Y�6���V�������T�}(r�EP螤  ���}H�E(   �]$�]r�M4Q��  ����^[��]�����U�����t]��]���������������̡����   ��ǀ�    V�p   �������������������������������U��E�� t��t3�]ù��"M �����]ø   ]����j j j jdjdhZ� j����?  � ����U���VWh`�jhjH�e�  ������t���R �N�(������3����H�A�U�R�Ћ��Q�Jj j��E�hL�P�у��U�R�M��X �8Vj�nB ��PWj j�`B ��PhZ� �BT ���M�����X ���H�A�U�R�Ѓ�_��^��]����������U��V��N蒹�����[Q �Et	V�Ϣ  ����^]� �����U���EV�����t	V訢  ����^]� ��������������U��U�BV�uW�}�g��'���F�g��'��������������AzT�M�B�f��&���A�f��&����������u.��!�B�a����!�G�a����������u_�   ^]� ��_3�^]� �������������U��M��t	��Pj��]������������U�����SV�U��Nh+Nd����*���������3�;ÉE�H���   �I����]��E�W�Vh��+Vd����*���������;�r�� �Nh+Nd�~d}�����*���������;�r�Y� �U��Fd�D�����G�U��C��;]���U��E��U�|�_���^[��]����������U��E��SV��Nh+NdW�}������*���������;�r�� �Fd�[�ЋU���M��Nh+ȸ���*���������;�r貾 �Vd�[�ʋM���Nh�E�+ʸ���*���������;�r聾 �Vd�E��[�D����`�U���M�� ���B�`�� �����^����z_^2�[��]� 3�9]~]�;]tQ;]tL;]tG�Nh+Nd�<�����*���������;�r�� �Vd��ʋM�U�P�E�QRP���A�����u��}C;]|�_^�[��]� ���������V��W���F|3�;�t	P藟  ���FpP�~|���   ���   �|�  �Fd��;�t	P�l�  ���NXQ�~d�~h�~l�W�  �FL��;�t	P�G�  ���V@R�~L�~P�~T�2�  ��_���^�������SVW��j���w@��  3ۃ�;�t�0�3���^�^�^j�wX��  ��;�t�0�3���^�^�^j�wp�Ŝ  ��;�t�0���_�^�^�^^[�3����_�^�^�^^[���������h�   膜  ����t���X���3�������U���S�ًKh+Kd����*����W��������]��y  3ɋǺ   ����V���Q�*�  ���ˋ��E� �J����P�����Au3���~'��$    ��@;�|��3���~�O���@I;�|��E����ߍ?�G���   ��M��E���I�M�����   ;؋ȉM�
�E�    �M�A;؉E�
�E�    �E��x;�3�VSWPQ�M��|�������   �}� �E�M������<��E�U�t-�M�E��E�P�����M�U��M��MR�����M�E��}�P�.�}��}�M�Q��������U�E�P�ωU�������M�U�M�R��������E�@;�}����L��@;�|�K��U�������V��  ��^_[��]� ��U��]�G����������U��M����w3ɍI���R蒚  ����]Ã��3����sލEP�M��E    �1� h���M�Q�E�x��~� �������U��E�U+���V�u��    +��~QRQV腸 ����^]�U��E�U+�V��W�}��    �49��vQRQW�S� ��_��^]� �����������U���E��P���\$�E�\$�E�$��]� �����������U��VW�����u赹 ���t��3ҋE�4@�G����;Bw��t�	�3�;As�� w��_^]� �������������U��E�U;�t.�MV�1�0�q�p�q�p�q�p�q�p�q�p��;�u�^]����U��M�U�E;�t.V�1�0�q�p�q�p�q�p�q�p�q�p����;�u�^]�U��U�M�E;�t0V�q���p�q���p�q�p�q�p�q�p�q�p;�u�^]���������������U��V��NP+NL����*��������W�}�;�r�m� �VL��ʍʋM�U��@_�^�@�E�]� ���������������U��V��NP+NL����*��������W�}�;�r�� �VL��ʍʋM�U��@_�^�@�E�]� ���������������U��E��t%�M���Q�P�Q�P�Q�P�Q�P�I�H]� �������������U����US�]V�uW�}2��E��M��E��E�PQRWVS����+󸫪�*��������@������ȋ�_^+�[��]�������U��j�h��d�    PQSVW�\�3�P�E�d�    �e��E�    �]�}�u��$    ;utVW���������}���u���E������ǋM�d�    Y_^[��]�j j �Ƕ ����������������U����US�]V�uW�}2��E��M��E��E�PQRWVS�R���+󸫪�*����������@��_^[��]����������������U��j�hЋd�    PQSVW�\�3�P�E�d�    �e��E�    �]�}�u��$    ��v�EPV��� ���O�}���u���E������M�d�    Y_^[��]�j j �ٵ ��U��Q�M�U�E� �E�P�EQ�MR�UPQR��������]�����U��Q�UV�uW�}�E� �E�P�ER��QPVW�)����v����_^��]� ��������U��SVW�}���    ��t�E9Fw;Fv�0� �E�]���G9^w;^v�� �]����t;�t� � �G;�t�VPRS�G������F��_^[]� ��������U��S�]V��W�    ��t�E9Fw;Fv谴 �E�}���C9~w;~v蔴 �}����t;�t耴 �S;�t/�F+�����    ���~QWQR蠲 ���E_�^^[]� _^��[]� ����������U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U���SV��FW�E�9Fv�� �~�;~v�ݳ �M��QSWP�U�R���r���_^[��]������������U���SV�ًCP�s@W�E�9Fv虳 �~��E�;~v至 �M��U�QRWP�E�P�������{h9{d�sXv�`� ��M�N�M�;Nv�K� �M��U�WRQP�E�P����������   9{|�spv�!� �^��M�;^v�� �U�WRSP�E�P���$���_^[��]��������������U��V�������Et	V蹔  ����^]� ���������������U��j�h��d�    P��$SVW�\�3�P�E�d�    �e���F��u3���V+и���*��������ȋ}���r  �^��+V����*��������º���
+�;�s������8;��  ���軪��
+�;�s�E�    �M��ȉM�;�s�U��j Q�0������ȉM�U+V����*����������E�    �EPW�[��P���'����E�   �MQ�UR�FP���m����E�   ߍ[�U��P�NQ�UR���K����E������^�N+˸���*������������t	S�?�  ���E�@�E�ȉV��ȉV�F�M�d�    Y_^[��]� �EP��  ��j j �� �ӋM+Ѹ���*���������;ǋE��   ��UЋP�UԋP�U؋P�U܋P�U��@�E�����E�PSQ���z����E�   �^�M�Q��+M����*���������+�WS��������E������EF�v�M�Q+�V�UR��������M�d�    Y_^[��]� ��MЋP�UԋH�M؋P�U܋H�M��P�U�<�����+ǉESSP��������FS�EP�MQ�6����U�R�E�WP�������M�d�    Y_^[��]� ���������������U���SV��^W�~��+ϸ���*���������u3��1;�v蒯 �M���t;�t耯 �M+ϸ���*����������M�U�EQjRP�������^;^v�H� �6W�M��u��]��p����E�M��U�_^��P[��]� ���������U���SV��^W��u3���N+˸���*��������ʋ~��+Ӹ���*���������;�s.�U�E� �M�Q�MR�FPQjW�l��������~_^[��]� ;�v蘮 �U�RWP�E�P������_^[��]� �����U����QP�E+QL��V�U��E�q@����*�����U��E���U��������u,���������Q�Y(�Q�Y0�Q �Y8�M�Q��� ���^��]� �������A������Au���Q���Q����z�Q�A ������Au���Q ���A(������z���Y(����A0������z���Y0����Q8����A�z����M���Q���{���^��]� ����U��E�E��$V3��0W���_�OP+OL����*�����������  S�OX�C����G(�g�G0�g�G8�g ��������Au.������Au%�؉u�������Au	�E   �o�   �E   �f������z2��������Au+���E�   ������Au3��E   �5�   �u�+����������E�   ����z3��E   ��u�   �OP+OL����*��OP+OL������򸫪�*���������u�d� �GL��vI�M�ȉU��U��؉M�А��E�M��]�� �U��]�R��OX�]������   EE�؃�u͋��   �wp�E9Fv��� �^��E�;^v�� �M�U�QRSP�EP�������V���F����N+N���������E��[�t�N+N����w衫 �F_^��]� _3�^��]� _��^��]� ��%��%��%��%���U��E��� ]��U����P�EP�EP�EPQ�J�у�]� �����������̡�V��H�QV�ҡ��H$�QDV�҃���^�����������U���V��H�QV�ҡ��H$�QDV�ҡ��U�H$�AdRV�Ѓ���^]� ��U���V��H�QV�ҡ��H$�QDV�ҡ��U�H$�ARV�Ѓ���^]� ��U���V��H�QV�ҡ��H$�QDV�ҡ��H$�U�ALVR�Ѓ���^]� �̡�V��H$�QHV�ҡ��H�QV�҃�^�������������U����P$�EPQ�JL�у�]� ����U����P$�R]�����������������U����P$�Rl]����������������̡��P$�Bp����̡��P$�BQ�Ѓ����������������U����P$��VWQ�J�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]� ���U����P$�EPQ�J�у�]� ����U����P$��VWQ�J �E�P�ы��u���B�HV�ы��B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�ҡ��H�A�U�R�Ѓ� _��^��]� ���U����P$��VWQ�J$�E�P�ы��u���B�HV�ы��B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�ҡ��H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e������Q$�JH�E�P�ы��B�P�M�Q�҃���^��]� ����̡��P$�B(Q��Yá��P$�BhQ��Y�U����P$�EPQ�J,�у�]� ����U����P$�EPQ�J0�у�]� ����U����P$�EPQ�J4�у�]� ����U����P$�EPQ�J8�у�]� ����U����UV��H$�ALVR�Ѓ���^]� ��������������U����H�QV�uV�ҡ��H$�QDV�ҡ��H$�U�ALVR�Ћ��E�Q$�J@PV�у���^]�U����UV��H$�A@RV�Ѓ���^]� ��������������U����P$�EPQ�J<�у�]� ����U����P$�EPQ�J<�у����@]� ���������������U����P$�EP�EPQ�JP�у�]� U����P$�EPQ�JT�у�]� ���̡��H$�QX�����U����H$�A\]�����������������U����P$�EP�EP�EPQ�J`�у�]� �����������̡��H(�������U����H(�AV�u�R�Ѓ��    ^]��������������U����P(�R]����������������̡��P(�B�����U����P(�R]�����������������U����P(�R]�����������������U����P(�R ]�����������������U����P(�E�RjP�EP��]� ��U����P(�E�R$P�EP�EP��]� ���P(�B(����̡��P(�B,����̡��P(�B0�����U����P(�R4]�����������������U����P(�RX]�����������������U����P(�R\]�����������������U����P(�R`]�����������������U����P(�Rd]�����������������U����P(�Rh]�����������������U����P(�Rl]�����������������U����P(�Rx]�����������������U����P(���   ]��������������U����P(�Rt]�����������������U����P(�Rp]�����������������U����P(�BpVW�}W���Ѕ�t:���Q(�Rp�GP���҅�t"���P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U����P(�BtVW�}W���Ѕ�t:���Q(�Rt�GP���҅�t"���P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U��VW�}W���0�����t8�GP���!�����t)�OQ��������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W���0�����t8�GP���!�����t)�O0Q��������t��HW��������t_�   ^]� _3�^]� ������������U������E�    �E�    �P(�RhV�E�P���҅���   �E���uG���H�A�U�R�Ћ��Q�E�RP�M�Q�ҡ��H�A�U�R�Ѓ��   ^��]� ���Qh�he  P���   �Ћ����E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�  ��3�^��]� �M��U�j IQ�MR������E�P��~  ���   ^��]� ���������������U�����V��H�A�U�R�Ѓ��M�Q������^��u���B�P�M�Q�҃�3���]� ���H$�E�I�U�RP�ы��B�P�M�Q�҃��   ��]� �U��Q���P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U����P(�R8]�����������������U����P(�R<]�����������������U����P(�R@]�����������������U����P(�RD]�����������������U����P(�RH]�����������������U����P(�E�R|P�EP��]� ����U����P(�RL]�����������������U����E�P(�BT���$��]� ���U����E�P(�BPQ�$��]� ����̡��H(�Q�����U����H(�AV�u�R�Ѓ��    ^]��������������U����P(���   ]��������������U����H(�A]����������������̡��H,�Q,����̡��P,�B4�����U����H,�A0V�u�R�Ѓ��    ^]�������������̡��P,�B8�����U����P,�R<��VW�E�P�ҋu�����H�QV�ҡ��H$�QDV�ҡ��H$�QLVW�ҡ��H$�AH�U�R�Ћ��Q�J�E�P�у�_��^��]� �������U����P,�E�R@��VWP�E�P�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� ��̡��H,�j j �҃��������������U����P,�EP�EPQ�J�у�]� U����H,�AV�u�R�Ѓ��    ^]�������������̡��P,�B����̡��P,�B����̡��P,�B����̡��P,�B ����̡��P,�B$����̡��P,�B(�����U����P,�R]�����������������U����P,�R��VW�E�P�ҋu�����H�QV�ҡ��H$�QDV�ҡ��H$�QLVW�ҡ��H$�AH�U�R�Ћ��Q�J�E�P�у�_��^��]� �������U����H��D  ]��������������U����H��H  ]��������������U����H��L  ]��������������U����H�I]�����������������U����H�A]�����������������U����H�I]�����������������U����H�A]�����������������U����H�I]�����������������U����H���  ]��������������U����H�A]�����������������U���V�u�E�P����������Q$�J�E�P�у���u-���B$�PH�M�Q�ҡ��H�A�U�R�Ѓ�3�^��]Ë��Q�J�E�jP�у���u=�U�R��������u-���H$�AH�U�R�Ћ��Q�J�E�P�у�3�^��]Ë��B�HjV�у���u���B�HV�у����I������Q$�JH�E�P�ы��B�P�M�Q�҃��   ^��]�����������U����H�A ]�����������������U����H�I(]�����������������U����H��  ]��������������U����H��   ]��������������U����H��  ]��������������U����H��  ]��������������U����H�A$��V�U�WR�Ћ��Q�u���BV�Ћ��Q$�BDV�Ћ��Q$�BLVW�Ћ��Q$�JH�E�P�ы��B�P�M�Q�҃�_��^��]������U����H���  ��V�U�WR�Ћ��Q�u���BV�Ћ��Q$�BDV�Ћ��Q$�BLVW�Ћ��Q$�JH�E�P�ы��B�P�M�Q�҃�_��^��]���U����H���  ]��������������U���<� SVW�E�    ��t�E�P�   �������/���Q�J�E�P�   �ы��B$�PD�M�Q�҃��}���H�u�QV�ҡ��H$�QDV�ҡ��H$�QLVW�҃���t)���H$�AH�U�R����Ћ��Q�J�E�P�у���t&���B$�PH�M�Q�ҡ��H�A�U�R�Ѓ�_��^[��]���U����H�U���  ��VWR�E�P�ы��u���B�HV�ы��B$�HDV�ы��B$�HLVW�ы��B$�PH�M�Q�ҡ��H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]����������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]�������������̡��H���   ��U����H���   V�uV�҃��    ^]�������������U����P�]����P�B����̡��P���   ��U����P�R`]�����������������U����P�Rd]�����������������U����P�Rh]�����������������U����P�Rl]�����������������U����P�Rp]�����������������U����P�Rt]�����������������U����P���   ]��������������U����P��  ]��������������U����P�Rx]�����������������U����P���   ]��������������U����P�R|]�����������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P�EPQ��  �у�]� �U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U��E��t ���R P�B$Q�Ѓ���t	�   ]� 3�]� U����P �E�RLQ�MPQ�҃�]� U��E��u]� ���R P�B(Q�Ѓ��   ]� ������U����P�R]�����������������U����P�R]�����������������U����P�R]�����������������U����P�R]�����������������U����P�R]�����������������U����P�R]�����������������U����P�E�R\P�EP��]� ����U����P�E��  P�EP��]� �U����E�P�B ���$��]� ���U����E�P�B$Q�$��]� �����U����E�P�B(���$��]� ���U����P�R,]�����������������U����P�R0]�����������������U����P�R4]�����������������U����P�R8]�����������������U����P�R<]�����������������U����P�R@]�����������������U����P�RD]�����������������U����P�RH]�����������������U����P�RL]�����������������U����P�RP]�����������������U����P���   ]��������������U����P�RT]�����������������U����P�EPQ��  �у�]� �U����P���   ]��������������U����P���   ]��������������U����P�RX]����������������̡��P���   ��U����P���   ]��������������U����P���   ]��������������U����P���   ]��������������U����P���   ]�������������̡��P���   ��U����P���   ]�������������̡��P���   ����P���   ����P���   ��U����H���   ]��������������U����H��   ]��������������U����H�U�E��VWRP���  �U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]������������U����H���  ]��������������U����P(�BPVW�}�Q�]���E�$�Ѕ�tM���G�Q(�]�E�BPQ���$�Ѕ�t,���G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U����P(�BTVW�}����$���Ѕ�tE���G�Q(�BT�����$�Ѕ�t(���G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U����P(�} �R8����P��]� �U����P�BdS�]VW��j ���Ћ��Q�����   h�Fh�  V�Ћ����E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ��Q(�BHV���Ѕ�t ���Q(�E�R VP���҅�t�   �3��EP�g  ��_��^[]� ������U���V�E���MP�k���P���#������Q�J���E�P�у���^��]� ��̡��P�BVj j����Ћ�^���������U����P�E�RVj P���ҋ�^]� U����P�E�RVPj����ҋ�^]� ���P�B�����U����P���   Vj ��Mj V�Ћ�^]� �����������U����P�EPQ�J�у�]� ����U����P�EPQ�J�у����@]� ���������������U����P�E�RtP�ҋ����   P�BX�Ѓ�]� ���U����P�E�Rlh#  P�EP��]� ���������������U����P�E�RlhF  P�EP��]� ���������������U����P�E�RtP�ҋ����   �M�R`QP�҃�]� ���������������U����P���   ]��������������U����P�E���   P�҅�u]� �����   P�B�Ѓ�]� ��������U���V�u�W�}�����Dz�F�_����D{:�F����$�:� �G��$�]��*� �E���������D{_�   ^��]�_3�^��]���������U���VW�M��`����E�}��t-���Q4P�B�Ѓ��M��u����_3�^��]Ë�R(����H0�QW�҃��M��tԋ�R Q�MQ���ҋ���P�B �M��Ѓ��t���Q0�Jx�E�PW�у��M��.���_��^��]�������U����P�B VW�}�����=NIVb��   ��   =TCAbtR=$'  t6=MicM��   ���Q���   j hIicM���ЋWP�B����_^]� ��BW����_�   ^]� ���Q���   j hdiem���ЋWP�B����_^]� =INIb��   �~ u���B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� �a�  _3�^]� =cnys����_3�^]� ������V���\����H0�Vh���҉F���F    ��^�����V��F�\���t���Q0P�B�Ѓ��F    ^�����̡��P0�A���   P�у����������U����P0�E�I���   PQ�҃�]� �������������̡��I�P0���   Q�Ѓ���������̡��P0�A���   j j j j j j j j j4P�у�(������̡��P0�A���   j j j j j j j j j;P�у�(�������U����P0�E�IPQ���   �у�]� ��������������U����E V��P�M��;������E�Q�R4Ph8kds�M��ҡ��E     �H0���   �U R�U�E�P�Ej R�UP�ER�UP�FRj2P�ыu ��(�M��������^��]� ��������������̡��I�P0���   Q�Ѓ����������U��V��F��u^]� ���Q0�M ���   j j j j j Q�Mj QjP�ҡ��H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uË��Q0P�B�Ѓ������̋A��u� ���Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5��v0Q�MQP���   R�U�R�Ћu�    �F    �����   j P�BV�Ћ����   �
�E�P�у�$��^��]� �������U����P0�E�I�RPQ�҃�]� �U��A��t)���Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5��v0QP���   R�Ѓ�^]� �����������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�V\�҃�^]� ����������U��A��u]� ���Q4�M��  Q�MQP�҃�]� �U��A��u]� ���Q4�M�RhQ�MQP�҃�]� ����U��A��u]� ���Q4�M�RpQ�MQP�҃�]� ����U��A��u]� ���Q4�M��  Q�MQP�҃�]� �U���$VW��htniv�M��I������P�E�R4Phulav�M��ҡ��P�B4hgnlfhtmrf�M��Ћ��E�Q�R4Phinim�M��ҡ��P�E�R4Phixam�M��ҡ��P�E�R4Phpets�M��ҡ��P�E�R4Phsirt�M��ҋE �}$=  �u�����t.���QP�B4h2nim�M��Ћ��Q�B4Wh2xam�M��ЋU�M�QR�E�P�����������   P�B8�Ћ����   �
���E�P�у��M��h���_��^��]�  ��������������U���$V��htlfv�M�������E���P�B,���$hulav�M��Ћ��E,�Q�R4Phtmrf�M����E���P�B,���$hinim�M����E���Q�B,���$hixam�M����E$���Q�B,���$hpets�M��Ћ��ED�Q�R4Phsirt�M��������E0��������Dzw���]8����Dzm�؋��E@�Q�R4Phdauq�M��ҋM�E�PQ�U�R���/��������   P�B8�Ћ����   �
���E�P�у��M�������^��]�@ �١��P�B,���$h2nim�M����E8���Q�B,���$h2xam�M����V�����U���$V��hgnrs�M��j����E���E��E�   �Q���   �E�Pj�M��ҡ����   ��U�R�ЋM���M����E�   �B���   �M�Qj�M��ҡ����   ��U�R�ЋU���M�QR�E�P�����������   P�B8�Ћ����   �
���E�P�у��M��������^��]� �U���$V��hmnrs�M��������P�E�R4Pj�M��ҋM�E�PQ�U�R�����������   P�B8�Ћ����   �
���E�P�у��M��n�����^��]� �����U��E��$�����VDSSS��P�M���������Q�B �M��Ћ��QjP�B4�M��ЋU�M�QR�E�P������������   P�B8�Ћ����   �
���E�P�у��M��������^��]� �����������U���$V��hCITb�M��j������P�E�R8PhCITb�M��ҡ��P�E�R4Phsirt�M��ҡ��P�E�R4Phulav�M��ҋM�E�PQ�U�R���<��������   P�B8�Ћ����   �
���E�P�у��M�������^��]� U��E��Vj ��P�M�Q�M������UPR���)�������H�A�U�R�Ѓ���^��]� ����������U��E,��UPj ���T$�$htemf�E$�� �\$�E�\$�E�\$�E�$R�/���]�( �����������U������E�������P��H���D{������������E��������D{����E,��Pj ���T$�U�$hrgdf�E$�� �������\$���\$�\$�E�$R����]�( ���������U��E,��Pj ���T$�U�$htcpf�E$�� �Ж�����\$�E���\$�}�\$�E�$R�C���]�( ���������������U��Q��u3�]� �E�E�H� V�5��v0Q�M Q�M���\$�E�$QPR�V(�҃�$^]� ������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�V,�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�V,�҃�^]� ����������U��Q��u3�]� �E�H� V�5��v0Q�MQPR�V0�҃�^]� ����������U��SVW���W��t$�E�H�5��^0� �uQVP�C0R�Ѓ���u	_^3�[]� �W��t��E�H� ���[0Q�NQPR�S0�҃���t̋W��tŋE�H� �=��0Q��VP�G0R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5��v0Q�MQ�MQPR�V<�҃�^]� ������U��QV3�W��u3��,�E�H� �5��v0Q�MQPR�V,��3Ƀ�9M��������M�B�P0VQ�M�ҋ�_^]� ����U��AV��u3��"�M�Q�	�5��v0R�URQP�F,�Ѓ������Q�E�M�R4PQ�M�ҋ�^]� ���������������U��A��V��u3��"�M�Q�	�5��v0R�U�RQP�F0�Ѓ������E��Q�E�M�R,���$P�ҋ�^��]� �����U�����V���U�V�U��]�W��t$�E�H� �=��0Q�M�QPR�W0�҃���u
_3�^��]� �V��t�E�H� �=��0Q�M�QPR�W0�҃���tˋV��tċE�H� �5��v0Q�M�QPR�V0�҃���t����P�M�RH�E�PQ�M��_�   ^��]� �����������U��� ��A�U�V�U�W�]���u3��&�M�Q�	�5��v0R�U�R�U�RQP�F<�Ѓ����E�}���t���Q�RH�M�QP���ҋE���t���E��Q���$P�B,����_��^��]� U����P�E���   Vj ��MP�ҋM$�U Q�MR�Uj Q�MR�UQPR������^]�  ����������U�����P�E���   V���$��MP���E8�E@�M,�Uj P���\$�E0�$Q�E$�� �\$���E�\$�E�\$�$R�����^]�< ������U�����P�E���   V���$��MP����Ej j ���T$���$htemf�E$�� �\$�E�\$�E�\$�$P����^]�$ �����������U�����P�E���   V���$��MP���E$�Ej �� �\$���E�\$�E�\$�$P����^]�$ ��������������U�����P�E���   V���$��MP����j j ���T$�E�$htcpf�E$�� �Ж�������\$�E���\$�}�\$�$P����^]�$ ���������������U����� V��H�A�U�R�ЋM�E��Qj �U�RP�M�Q�M��h���UPR�����������H�A�U�R�Ћ��Q�J�E�P�у���^��]� ������������U���dV��M��������Q���   P�EP�M�Q�M��P�M������M��Q���j j �E�P�M������MPQ���U��������B�P�M�Q�҃��M������M�������^��]� �����U���P��EV�]���W�}����t���Q���$P���   �����]�����U��UЍE��]؋Q�M���   PQ�E�P���ҋ�M��P�U�H�M�P�U�H�M��P�F�U��u_^��]� �M�E�Q�	�5��v0R�U R���\$�U��E��$RQP�F(�Ѓ�$_^��]� ���������������U���0�E�M���u���H���   �҅�u��]� SVW���_  ��htlfv�MЉu�z����E�}���X�U�����$�̂ �]��G�$辂 �}�S,�M��$hulav�ҡ��P�B4hmrffhtmrf�M��Ћ}����M�Y���$�u� �]��G�$�g� �}�S,�M��$hinim�ҋ}����M�X���$�9� �]��G�$�+� �}�S,�M��$hixam������P�B,���$hpets�M��Ћ��Q�B4j hdauq�M��Ћ��Q�B4Vhspff�M��Ћ��E �Q�R4Phsirt�M��ҋM�E�PQ�M��U�R�^��������   P�B8�Ћ����   �
���E�P�у��M��;���_��^[��]� U��E��V���u���H���   �҅�u^��]� ���N]  �E�F��u3��"�M�Q�	�5��v0R�U�RQP�F0�Ѓ����E������M������\$�M��$�
 ��M��P�Q�P�Q�@�A��^��]� ����������U���0����]�V���M�]�P���   �E�PQ�M�E�P�ҋ�P�M��Hj �U�P�E P�M��MQ�M�U��UR�U�E�PQR������^��]� ���������������U�����UV�]���E�P�]��ERP�������Q�M�R@���E�PQ�M�ҋ�^��]� ����������U��A��u]� �M�Q�	V�5��v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� ���Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� ���Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U����P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� ���Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj>P�ҋE���(��]� ������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5��v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M�� �MQ�U�R�M��� ��tm�}��E��tN�����   P�BH�ЋM��I����tQ�W�7���[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M��{ ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5��v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� ���E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� ���Q0�M�RDQ�MQ�MQP�҃�]� U��A��u]� ���Q0�M�RHQ�MQ�MQ�MQ�MQ�MQP�҃�]� ���̋A��uË��Q0P�BX�Ѓ�������U��A��u]� ���Q0�M�RLQ�MQP�҃�]� ����U��A��u]� ���Q0�M�RP��   �QP�҃�]� ��U��A��u]� ���Q0�M�RPQP�҃�]� ��������U��A��u]� ���Q0�M�RTQ�MQ�MQ�MQP�҃�]� ������������U���V�u�VW���H4�R�ЋE�F    �~�H� ���R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� ���Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I���R0P�EPQ���   �у�]� ������̡��I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u��� ���R0�I�R@V�uVP�EPQ�҃�^]� �����������U����P0�E�I�RdP�EP�EP�EP�EPQ�҃�]� �U����P0�E�I�RpP�EP�EP�EP�EPQ�҃�]� �U��E�P� V�5��v0R�UR�UR�UR�URP�A�NhP�у�^]� ��������U��E� ���R0j j j j j j j P�A���   jP�у�(]� �����������U��E� ���R0j j j j j jj P�A���   jP�у�(]� �����������U��E� ���R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M������E�H� ���R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R������M�������^��]� ����������U��E�P� V�5��v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5��v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5��v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5��v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U����P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U����UVj j j j j R��H0�E�Vj P���   jR�Ћ��Q0�E�N�RtPQ�҃�0^]� ��U����P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡��P0�A���   j j j j j j j j jP�у�(�������U����P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡��P0�A���   j j j j j j j j j(P�у�(�������U����P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U����P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡��P0�A���   j j j j j j j j jP�у�(������̡��P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}�M���t���P���   j j���Љ�u��t���Q���   j j���Љ���Q0�E��H�R`VWQ�҃�_^[��]� �U����P0�E�I���   P�EP�EPQ�҃�]� �����̡��P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V���\����H0�Vh���҉F3��F�F������F   ��^�������V��F�\���t���Q0P�B�Ѓ��F    ^������U��E�UVj ��MP�EQ3�9MR��Pj �F    ��
Q��������t�~ t
�   ^]� 3�^]� �U��E�A�I��u3�]� ���B0Q�H�у�]� ����U����P�B S�]V�����=ckhc��   ��   =cksate=TCAb��   ���Q���   Wj hdiem���Ћ���BSW���F   �Ѓ~ ��t��t��u3Ƀ���Q���C���_^��[]� �~ tK��B����^[]� �~ t6��������t+�F    ^�   []� =atnit�MQS������^[]� ^3�[]� �U��V��~ ��   W�}����   �$���E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN���M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W��d  ���F    _^]� D�R�`�n�|�������������U��V��~ �  �E W�}�E����   �$�p����]������   �   ���]����A��   �   ���]����A��   �r���]������   �`�E������A��uN��������   �C�E��������u1������A{{�*�E���������E������A�����]����DzU����ء��U�H0�F���   j j j j j j j RjP���E �U(��(R���\$�E�$W�c  ���F    _^]�$ �I j���������������������������U���E �E�Uj���\$�E�\$�E�$PR�w���]�  ���U���E �E�Uj���\$�E�\$�E�$PR�G���]�  ���U���E �E�Uj���\$�E�\$�E�$PR����]�  ��̋�3�� Ĝ�H�H�H�������������VW��3��Ĝ9~u���H4�V�R�Ѓ��~�~_^����U����P4�E�I�RtPQ�҃�]� �U��U��t3�A���I0R���   P�ҋ��Q0�M���   QP�҃�]� ���P0�E�I�R|PQ�҃�]� ������̡��P4�A�JP�у������������̡��P4�A�JP�у������������̡��P4�A�JP�у������������̡��P4�A�J|P�у������������̡��P4�A���   P�у����������U����P4�E�I�RP�EP�EP�EPQ�҃�]� �����U����P4�E�I�RP�EP�EP�EPQ�҃�]� �����U����P4�E�I�R PQ�҃�]� �U����P4�E�I�R$PQ�҃�]� �U����P0�E�I���   P�EP�EP�EPQ�҃�]� ��U����P4�E�I���   PQ�҃�]� ��������������U����P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U����P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U����P4�E�I�R(PQ�҃�]� �U����P4�E�I�R,P�EP�EPQ�҃�]� ���������U����P4�E�I�R0P�EPQ�҃�]� ������������̡��P4�A�J4P��Y��������������U����UV��EP�M�Q�NR�E�    �E�    �������H4�V�AR�Ћ��Q0�Rhj �M�Q�M�Q�M�Q�M�QP�F�HQ�҃� �} ^t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ��������������U����P4�E�I�R8PQ�҃�]� �U����P4�E�I�R<PQ�҃�]� �U����P4�E�I���   P�EPQ�҃�]� ����������U����E�P4�A��  ���$P�у�]� ��������̡��P4�A�J@P�у������������̡��P4�A��  P�у����������U����P4�E�I�RDP�EPQ�҃�]� �������������U����P4�E�I�RHP�EPQ�҃�]� �������������U����P4�E�I�RLP�EPQ�҃�]� �������������U����P4�E�I�RPP�EPQ�҃�]� �������������U���SV�uW�����   �QV�҃�����   �����   �]�QS�҃�S��uA�����   �Q@�ҋء����   �Q@V�ҋ��Q4�JPSP�GP�у�_^[]� �����   �H�у���uD�����   �H8S�ы��؋��   �H@V�ы��J4�WSP�AHR�Ѓ�_^[]� h�h�  ��   �����   �BV�Ѓ�����   �����   �]�BS�Ѓ�S��uC�����   �B@�Ћ����   �؋B8V�Ћ��Q4�JLSP�GP�у�_^[]� �����   �H�у���uD�����   �H8S�ы��؋��   �H8V�ы��J4�WSP�ADR�Ѓ�_^[]� h�h�  �
h�h�  ���Q��0  �Ѓ�_^[]� �U����P4�E�I��  P�EP�EP�EPQ�҃�]� ��U����P4�E,P�E(P�E$P�E �IP�E�RTP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U����P4�E�I�RXP�EP�EP�EPQ�҃�]� ����̡��P4�A�J`P��Y�������������̡��P4�A�JdP�у�������������U����P4�E�I��   P�EP�EP�EPQ�҃�]� ��U����P4�E�I�R\P�EP�EP�EP�EP�EPQ�҃�]� �������������U����P4�E�I�RhP�EPQ�҃�]� �������������U����P4�E�I��  P�EPQ�҃�]� ����������U����P4�E�I��  P�EPQ�҃�]� ����������U����P4�E�I�RpP�EPQ�҃�]� �������������U���,V��~ ��   ���V�H4�AR�Ѓ} t ���Q0�RlP�F�HQ�҃�^��]� ��hARDb�MԉE��E�    �\���P�M�Q�N�U�R�{��������   ��U�R�Ѓ��M��m���^��]� ������U����P4�E�I�RlPQ�҃��   ]� ������������U����E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U����P4�E�I���   P�EP�EPQ�҃�]� �����̡��P4�A���   P�у���������̸   ����������̸   �����������U���V��H4�V�A$h�  R�Ћ��Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U����P4�E�I�RxP�EP�EP�EPQ�҃�]� �����U����P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}�M���t���P���   j j���Љ�u��t���Q���   j j���Љ���Q4�E��H�RpVWQ�҃�_^[��]� �U��Q���P�B SVW�}���3���=INIb�/  �  =SACbvt+=$'  t
=MicM�  ��B$W����_�   ^��[��]� ��R3��E��E�EP�M�Q���҅�t���U�H4�E�R�VP�AR�Ѓ�_�   ^��[��]� =ARDb�  ���Q���   j j���Ћ��Qj �؋��   j���Ћ��Qj �E����   j���Ћ��Qj �E���   j���ЋM���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>���I���P���!���P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� ���Q���   j hIicM���ЋWP�B ����_^[��]� �������������U����P4�E�I�RTh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M��:������Q4�JlP�FP�у��M��\���^��]��������V���\����H0�Vh���҉F���F    �4��F   ��^��������V��F�\���t���Q0P�B�Ѓ��F    ^������U����P�B VW�}�����=cksat`=ckhct�MQW��荽��_^]� �Nj j j j j j �F   ���B0���   j j j Q�҃�(��t'_�F    �   ^]� �~ t��P����_^]� _3�^]� ���U����H���  ]��������������U����H0���   ]��������������U����H0�U�E��VWRP���   �U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]������������U����H0���   ]��������������U����H0���   ]��������������U����H0���   ]��������������U��Ej0P�K  ��]��������������U��Ej0P�r�  ��P�iK  ��]�����U��E�M��j0PQ�U�R�w�  ��P�>K  ���H�A�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P��  ��P��J  ���Q�J�E�P�у���]��U��Ej$P��J  3Ƀ�������]����U��Ej$P��  ��P�J  3Ƀ�������]�����������U��E�M��Vj$PQ�U�R��  ��P�mJ  ��3Ƀ��B�P����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P���  ��P�J  ��3Ƀ��B�P����M�Q�҃���^��]����U����H�U�E���   RPj �у�]���������������U����H�U�ER�UP���   Rj �Ѓ�]�����������U����P4�E�I�R,P�EP�EPQ�҃�]� ���������U����P4�E�I�R0P�EPQ�҃�]� ������������̡��P4�A�J4P��Y��������������U��U��V��EP�M�QR���4������H0�E�P� R�U�R�U�R�U�R�U�R�VP�AhR�Ѓ��} ^t(�} t(�E�M�;�~<�U��;�}3�E�M�;�~)�U���} u�E�M�;�~�U��;�}�   ��]� 3���]� �����������U��ESVW�؅�u�Y���P�}���   j hdiuM���Ћ���tK;3u	_^3�[]� ���Q���   j hIicM����;�u���Q���   j h1icM���Шu��3_^�   []� �����U����P�BT��(V�uhfnic���Ѕ�t���Q�ȋ��   j
�Ѕ���   ���Q�RPhfnic�E�P����P�M��ߴ���M�������u�E�P��������M��������Q�B ���Ѓ��t���Q�B ���Ѕ�u���Q�B$hfnic���Ћ��E�Q�R8Pj
����^��]���������U����P0�E�IP�EP�EP�EPQ���   �у�]� ��U����P0�E�IV�p� ���   V�uj j j V�uVj Pj=Q�҃�(^]� ����U����P0�E�IV�p� ���   V�uV�uj j j�Vj Pj=Q�҃�(^]� ���̡��I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V���\����H0�WVh���ҋ}�F�E�F    �F   �\��F���Q���   ��j hmyal���ЉF��t��t�F    ���Q���   j
hhfed���ЉF_��^]� �����������U����P�B VW�}�����=ytsdt�MQW�������_^]� ���B0�N���   Q�ҋ�P������_�   ^]� ��3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ��������������������̸�������������U���E�Y(]� ���U���(V���P(�M�Q���ҋN��t&���R0j j j j j j P���   j jQ�Ѓ�(���Q�J�E�P�ы��B�P�M�Q�ҋF����t ���Q0�RHj �M�Qj jj?j P�҃����H�A�U�WR�Ћ��Q�J�E�P�ыF����u3��;���E�    �J0�U�Rj j j h  
 j�U�Rh�  jP���   �Ћ}���(���Q�J�E�P�у���_u3�^��]Ë��B�P�M�Q�ҋF����t ���Q0�RHj �M�Qj j j8j P�҃����H�A�U�R�ЋF����t���Q0jP�BP�Ѓ����Q�J�E�P�у��M�詯��Ph   h  K j;�U�Rh	��h�  ���w������H�A�U�R�Ѓ��M��˯���F��t���Q0P�BX�Ѓ��F��t���Q0P�BX�Ѓ��F��t'���Q0j j j j j jj j jP���   �Ѓ�(j�v$�QA  ���   ^��]�����U���SV��W�~j����  ��V�^(3ۉ^4�^8�^<���H0�Ah�   R�Ћ��Q�J�E�P�ы��B�PSj��M�h��Q�҃�SS�E�P�M�Q���E��  �]��	������B�P�M�Q�҃�Sj�����  _^[��]���̍A�������������U��VW��~4 tA�I ���H��0  h�hs  ��j
�oJ  ���HP�V �AR�Ѓ���uQ9F4u��QP�Bh�~0���Ѓ~4 t;���Q��0  h�h�  �Ћ��QP�Bl�������m���_3�^]� �M�U�N8�V4���PP�Bl�~0���Ѓ~4 t%j
��I  ���QP�F �JP�у���u�9F4uۋ��BP�PhS���ҋ^<�F<    ���PP�Bl���Ћ�[_^]� ��U����P�B ��@VW�}�����=MicMtI=fnic��   j�M�������uP���=����M��%������Q�B4jj����_�   ^��]� ���Q���   j hIicM����=�����   htats�M�蒬�����Q�B0j j�M��ЍM�Q�U�R�E�P���E��  �E�    茳�������   �
�E�P�у��M��}����F�F   ��t���J0�QP�҃��EPW���1���_^��]� ���������U��E��V��t3�^]� j�N��  j�
>  �F    �v����t���H0�QV�҃��   ^]� ��������������j���V�  j�=  ��3�����������U��E3�h�����h  ���P�Ej BR�Uj PR�����]� �U��Q�Q��u3���]� �E�H� V�5�Q�M�Q�E�    �v0PR�V8�ҋ�����t@�E���t9���Q�M�RQP�ҋE�����t���QW��P�B��W�S  ��_��^��]� ������U�����V��H�A�U�R�ЋU���M�QR���D�������u���H�A�U�R�Ѓ�3�^��]� �M�Q�M�������B�P�M�Q�҃���^��]� �������U�����V��H�A�U�R�ЋU���M�QR��������M����P�R8�E�PQ�M�ҡ��H�A�U�R�Ѓ���^��]� �������������U���V��M��/����M�E�PQ������������B�U�@<�M�Q�MR�ЍM�������^��]� ����U����P�E���   Vj ��MP��h���h  �j j jj P�EP������^]� ��������������U���V�uW�����   �QV�҃�V��u,�����   �Q@�ҋ��Q4�J P�GP�у�_^]� �����   �H�у���u.�����   �H8V�ы��J4�WP�A$R�Ѓ�_^]� ���Q��0  h�h  �Ѓ�_^]� �����U���4���H�QSVW�}W�ҡ��P�u���   ��3�SS�Ή]�Ћ��QS�E����   j���Ћ�;��L  �d$ �} ~l���Q�J�E�P�ы��B�Pj j��M�hĝQ�ҡ��P�B<�����Ћ��Q�RLj�j��M�QP���ҡ��H�A�U�R�Ѓ����Q0�E����   VP�M�Q�ҋ���H�A�U�R�Ћ��Q�J�E�PV�ы��B�P�M�Q�ҡ��P�B<�����Ћ��Q�RLj�j��M�QP���ҡ��H�A�U�R�Ћ��Q�u���   �E��j ��
S���Ћ��Q���   �E�j �CP���ҋ����������_^[��]����������������U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj AQj R�UR������^]� ��������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR�ϯ��^]� ����������U��E�E43҃8��R�U<R�U(���\$�E,�$R�E �� �\$�E�\$�E�\$�@�E�$P�°��]�8 ��������������U��E�@3҃8��E��Rj ���T$�$htemf�E �� �\$�E�\$�E�\$�$P�g���]�  ���U��E�E 3҃8��R�� �\$�E�\$�E�\$�@�E�$P�
���]�  ������U��E�@3҃8��E��Rj ���T$�$htcpf�E �� �Ж�����\$�E���\$�}�\$�$P�˯��]�  �������U��E3҃8��R�UR�UR�UR�UP�EPR����]� U��E3҃8V�u��V��RP�EP�����^]� ����������U��Q��u3�]� �E�E�H� V�5��v0Q�M Q�M���\$���E�$QPR�V(�҃�$^]� ���U����P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U����P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U�����P�E���   V���$��MP�ҋ���u�^�    ^]� ��u�^����D{�   ^]� ��^]� ������U���0����U�V�U���M�]��P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�Q�P�Q�P�@�Q�A����  ^��]� ��������U��� ����]�V���M�]��P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�@�Q�A����  ^��]� �����U���VW�}�M�;}us���P�u���   j htsem���Ѕ�uS���QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E��������t�E�M�P�w  _�   ^��]� _3�^��]� U���VW�}�M�;}us���P�u���   j htsem���Ѕ�uS���QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E�跲����t�E�M�P��  _�   ^��]� _3�^��]� U���SVW�}��;}uz���P�u���   j htsem���Ѕ�uZ���QP���   hrdem���Ѕ�u=��M�Q�]��M�U�R�}��E��e�����t�E������$�  _^�   [��]� _^3�[��]� ��������U���4�ESW�}�M�;�t;Et	;E��   ���P�]���   j htsem���Ѕ���   ���QP���   hrdem���Ѕ�uj�M��U�ỦE��UԉE��]܉E�M�E�P�M�Q�M�U�U�R�E�P�}��ѱ����t+�E̋M�������E��X�E��X��  �   _[��]� _3�[��]� ��������U���SVW�}��;}��   ���P�u���   j htsem���Ѕ�uj���QP���   hrdem���Ѕ�uM��U�M��]���Q�M�]��E�R�E�P�}��H�����t%�E��������E��X�  �   _^[��]� _^3�[��]� ���̋A���X(Q�ȋB$��j j h���� 4  ���������������U�����0VW���H�A�U�R�Ћ��Q�J�E�P�ыE���U�RP�M�Q�M�������J�U�RP�A�Ћ��Q�J�E�P�ы��B�P�M�Q�ҡ��H�Q��V�ҡ��H�A�U�VR�Ѓ�����  ���Q�J�E�P�у�_^��]� ������������U���SVW�}��;}��   ���P�u���   j htsem���Ѕ�ue���QP���   hrdem���Ѕ�uH���Q�J�E�P�ыM���U�R�E�P�}��E�    �-�����u ���Q�J�E�P�у�3�_^[��]� ���U��R�;�����  ���H�A�U�R�Ѓ�_^�   [��]� ��U��V�u���  ��^]� �����������U���L��SV��H�A�U�R�Ћ��Q�J3�Sj��E�hȝP���F(�Ж��S�U�SR�E��  �]��H: P�E�P�n1����P�M�Q�Q�����P�U�R���������H�A�U�R�Ћ��Q�J�E�P�ы��B�P�M�Q�҃�htats�M��=������P�B0jj�M����F(���Q�B,���$j�M��ЍM�Q�U�R�E�P���E��  �]�� ��������   �
�E�P�у�9^4t^���BP�PhW�~0���ҋF4;�t�N8Q�Ѓ��F<�^8�^4����B��0  h�h�  �у����BP�Pl����_�M�讛��^[��]� ������U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�E�Y����D{�   ]� �����������U�����u�E�    �Y�E�Y�E�Y]� ��u-�E�Y����Dz�E�Y����Dz�E�Y����D{�   ]� �����U��V�����u#�E�M�U�F�E�N�V�    �F^]� ��u�MQ�VR�O�������t�   ^]� �������������U��V��~ �Ĝu���H4�V�R�Ѓ��E�F    �F    t	V�q  ����^]� �������U��V��F�\���t���Q0P�B�Ѓ��E�F    t	V�(  ����^]� ��������������U���V��3ɍF��H��������M��M����   �RQ�M�QP�ҡ����   ��U�R�Ѓ���^��]��������������U��V�����u �    ���H�A���UVR�Ѓ��#��u���Q�Rx�EP�N�҅�t�   ���H�A�UR�Ѓ�^]� �������U��V�u���t���QP��Ѓ��    ^]���������̡��H��@  hﾭ���Y����������U��E��t���QP��@  �Ѓ�]����������������U����H���  ]��������������U����H��  ]�������������̡��H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�R6 ������u_^]Ã} tWj V�, ��_������F��   ^]���U����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW��5 ������u_^]�Wj V� ��_������F��   ^]�������������U����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�V5 ������u_^]�Wj V�6 ��_������F��   ^]�������������U����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW��4 ������u_^]�Wj V� ��_������F��   ^]�������������U����E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�V4 ������u_^]�Wj V�6 ��_������F��   ^]�������������U��M��t-�=� t�y���A�uP�Q ��]á��P�Q�Ѓ�]��������U��M��t-�=� t�y���A�uP� ��]á��P�Q�Ѓ�]��������U����H�U�R�Ѓ�]���������U����H�U�R�Ѓ�]���������U����E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�3 ������u_^]�Wj V�� ��_������F��   ^]���������U����E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   ����t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�#2 ������u_^]�Wj V� ��_������F��   ^]����������U��E��w�   ����t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�1 ������u_^]�Wj V�p ��_������F��   ^]�������U����H�U�R�Ѓ�]���������U����H�U�R�Ѓ�]���������U����H�U�R�Ѓ�]���������U����H�U�R�Ѓ�]��������̡��HL���   ��U����H@�AV�u�R�Ѓ��    ^]�������������̡��HL�������U����H@�AV�u�R�Ѓ��    ^]�������������̡��PL���   Q�Ѓ�������������U����PL�EP�EPQ���   �у�]� �������������U���V��HL���   V�҃���u���U�HL���   j RV�Ѓ�^]� �����   �ȋBP�Ћ����   �MP�BH��^]� �����̡��PL��(  Q�Ѓ�������������U����PL�EP�EPQ��,  �у�]� ������������̡��HL�Q�����U����H@�AV�u�R�Ѓ��    ^]��������������U����PL�E�R��VPQ�M�Q�ҋu��P���e����M��}�����^��]� ����U����PL�EPQ���   �у�]� �U����PL�EP�EPQ�J�у�]� ���PL�BQ�Ѓ���������������̡��PL�BQ�Ѓ���������������̡��PL�BQ�Ѓ����������������U����PL�EP�EP�EPQ�J �у�]� ������������U����PL�EPQ��4  �у�]� �U����PL�EP�EP�EPQ�J$�у�]� ������������U����PL�EP�EP�EP�EPQ�J(�у�]� �������̡��PL�B,Q�Ѓ���������������̡��PL�B0Q�Ѓ����������������U����PL�EP�EPQ��  �у�]� ������������̡��PL���   Q�Ѓ�������������U����PL�E��  ��VPQ�M�Q�ҋu��P���B����M��Z�����^��]� ̡��PL�B4Q�Ѓ���������������̡��PL�B8j Q�Ѓ��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL��l  ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL���   ]��������������U����PL�EPQ�J<�у�]� ���̡��PL�BQ��Y�U����PL�EP�EPQ�J@�у�]� U����PL�Ej PQ�JD�у�]� ��U����PL�Ej PQ�JH�у�]� ��U����PL�EjPQ�JD�у�]� ��U����PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��E  W�M�Q�U�R���tM  ���M����7  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  ��D  j�M�Q�U�R����L  �M���6  �����   ��U�R�Ѓ�^��]�����������U���$���UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��zD  j�E�P�M�Q���YL  �M��q6  �����   ��M�Q�҃�_^��]� ��U���$���UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}���C  j�E�P�M�Q����K  �M���5  �����   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��C  W�M�Q�U�R���TK  ���M����5  ��t+�u���f�������   ��U�R�Ѓ�_��^[��]� �����   �JL�E�P�ыu��P���%g�������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}���B  W�M�Q�U�R���J  ���M�����4  ��t+�u����e�������   ��U�R�Ѓ�_��^[��]� �����   �JL�E�P�ыu��P���ef�������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��B  W�M�Q�U�R����I  ���M����4  _^��[t�����   ��U�R�������]Ë����   �J<�E�P���]������   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��dA  W�M�Q�U�R���$I  ���M����W3  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��@  W�M�Q�U�R���tH  ���M����2  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� �����̡��PL���   Q��Y��������������U����PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U����PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��$?  W�M�Q�U�R����F  ���M����1  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��T>  W�M�Q�U�R���F  ���M����G0  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��=  W�M�Q�U�R���DE  ���M����w/  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��<  W�M�Q�U�R���tD  ���M����.  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  ��;  j�M�Q�UR����C  �M��-  �����   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��;  j�U�R�E�P���nC  �M��-  �����   �
�E�P�у�^��]� ��������U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
;  j�E�P�M�Q����B  �M��-  �����   ��M�Q�҃�_^��]� ��U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��:  j�E�P�M�Q���iB  �M��,  �����   ��M�Q�҃�_^��]� ��U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
:  j�E�P�M�Q����A  �M��,  �����   ��M�Q�҃�_^��]� ��U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��9  j�E�P�M�Q���iA  �M��+  �����   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��9  j�U�R�E�P����@  �M��+  �����   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}��8  W�M�Q�U�R���t@  ���M����*  ��t-��u������   ���^�U�R�Ѓ�_��^[��]� �����   �JP�E�P�ы�u�H��P�@�N���V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���7  W�M�Q�U�R���?  ���M�����)  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��47  W�M�Q�U�R����>  ���M����')  ��t�����   ��U�R�Ѓ�_^3�[��]Ë����   �J8�E�P�ы������   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ���̡��PL���  ��U���$���UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��:6  j�E�P�M�Q���>  �M��1(  �����   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���5  j�U�R�E�P���=  �M���'  �����   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��_5  j�U�R�E�P���>=  �M��V'  �����   �
�E�P�у�^��]� ��������U����H���   ]��������������U����H���   ]�������������̡��H���   ����H���   ��U����H���   V�u�R�Ѓ��    ^]�����������U����H���   ]��������������U����HL�QV�ҋ���u^]á��H�U�Ej R�UP��h  RV�Ѓ���u���Q@�BV�Ѓ�3���^]��������U����H�U�E��h  j R�U�� P�ERP�у�]����U����H���   ]��������������U����H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡��PL�BLQ�Ѓ���������������̡��PL�BPQ�Ѓ����������������U����PL�EP�EPQ�JT�у�]� U����PL�EPQ��  �у�]� �U����PL�EPQ���   �у�]� ̡��PL�BXQ�Ѓ����������������U����PL�EP�EP�EPQ�J\�у�]� ������������U���4��SV��HL�QW�ҋ�3ۉ}�;��x  �M��!x�����E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ����   �BSSW���Ѕ���   ���QL�BW�Ћ���;���   ��    �����   �B(���ЍM�Qh�   ���u��j  ������   �M�;���   �����   ���   S��;�tm�����   �ȋB<V�Ћ����   ���   �E�P�у�;�t���B@�HV�у���;��\����}��M��!  �M��Yw����_^[��]� �}����B@�HW�ы����   ���   �M�Q�҃��M��9!  �M��w��_^3�[��]� �����̡��PL�B`Q�Ѓ���������������̡��PL�BdQ�Ѓ����������������U����PL�EPQ�Jh�у�]� ���̡��PL��D  Q�Ѓ������������̡��PL�BlQ�Ѓ����������������U����PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh`h@h hR�Q�U R�UR�UR�U���A�$�5��vLRP���   Q�Ѓ�4^]�  ������̡��PL���   Q�Ѓ�������������U����PL�EP�EP�EPQ��   �у�]� ���������U����PL��H  ]�������������̡��PL��L  ��U����PL��P  ]��������������U����PL��T  ]��������������U����PL��p  ]��������������U����PL��t  ]��������������U����PL�EP�EP�EP�EP�EPQ���   �у�]� �U����PL�EP�EP�EPQ���   �у�]� ���������U����PL�EP�EP�EP�EPQ��   �у�]� �����U����HL���   ]��������������U����HL���   ]��������������U����HL���   ]�������������̡��HL��  ����HL��@  ��U����PL���  ]��������������U����PL���  ]��������������U����PL���  ]��������������U��� ��V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\���QLjP���   ���ЋM��U�Rh=���M�}��  �������   ���   �U�R�Ѓ��M��u��  ��_^��]Ë����   ���   �E�P�у��M��u��^  _�   ^��]����U��� ��V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\���QLjP���   ���ЋM��U�Rh<���M�}��C  �������   ���   �U�R�Ѓ��M��u��  ��_^��]Ë����   ���   �E�P�у��M��u��  _�   ^��]����U����P8�EPQ�JD�у�]� ���̡��H8�Q<�����U����H8�A@V�u�R�Ѓ��    ^]�������������̡��H8�������U����H8�AV�u�R�Ѓ��    ^]��������������U����P8�EP�EP�EPQ�J�у�]� ������������U����P8�EP�EPQ�J�у�]� ���P8�BQ�Ѓ����������������U����P8�EPQ�J �у�]� ����U����P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U����P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U����P8�EP�EPQ�J(�у�]� U����P8�EP�EP�EPQ�J,�у�]� ������������U����P8�EP�EP�EPQ�J�у�]� ������������U����P8�EP�EP�EP�EP�EPQ�J�у�]� ����U����P8�EP�EPQ�J0�у�]� U����P8�EP�EP�EPQ�J4�у�]� ������������U����P8�EPQ�J8�у�]� ����U����H��x  ]��������������U����H��|  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H�A,]�����������������U����H���  ]��������������U����H�QV�uV�ҡ��H�Q8V�҃���^]�����̡��H�Q<�����U����H�I@]����������������̡��H�QD����̡��H�QH�����U����H�AL]�����������������U����H�IP]�����������������U����H��<  ]��������������U����H��,  ]��������������U����H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡��H���   ����H���  ��U����H�U�ER�UP�ER�UP���   Rh�2  �Ѓ�]����������������U����H�A]�����������������U����H��\  ]��������������U����H�AT]�����������������U����H�AX]�����������������U����H�A\]����������������̡��H�Q`�����U����H���  ]�������������̡��H�Qd����̡��H�Qh�����U����H�Al]�����������������U����H�Ap]�����������������U����H�At]�����������������U����H��D  ]��������������U����H��  ]��������������U����H�Ix]�����������������U����H��@  ]��������������U��V�u���G�����H�U�A|VR�Ѓ���^]���������U����H���   ]��������������U����H��h  ]��������������U����H��d  ]��������������U����H���  ]�������������̡��H���   ��U����H��l  ]��������������U����H��   ]��������������U����H��  ]��������������U��V�u����h�����H���   V�҃���^]���������̡��H��`  ��U����H��  ]��������������U����H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U����H���  ]��������������U��U�E���H�E���   R���\$�E�$P�у�]�U����H���   ]��������������U����H���   ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���   ]��������������U����H���   ]��������������U����H���   ]��������������U����H���   ]��������������U����H���   ]��������������U����H���   ]��������������U����P���E�P�E�P�E�PQ���   �у����#E���]����������������U����P���E�P�E�P�E�PQ���   �у����#E���]����������������U����P���E�P�E�P�E�PQ���   �у����#E���]����������������U����H��8  ]��������������U��V�u(V�u$�E�@���R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@���R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U����P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U����P0�EP�EP�EP�EPQ���   �у�]� ����̡��P0���   Q�Ѓ�������������U����P0�EP�EPQ���   �у�]� �������������U����P0�EP�EP�EP�EPQ���   �у�]� ����̡��P0���   Q�Ѓ������������̡��H0���   ��U����H0���   V�u�R�Ѓ��    ^]�����������U����H��H  ]��������������U����H��T  ]�������������̡��H��p  ����H���  ��U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H�U�E��X  ��VR�UPR�E�P�ыu�    �F    �����   �Qj PV�ҡ����   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M��Jb��P�E�hicMCP�k������M��pb�������   �JT�E�P�у���u(�u����a�������   ��M�Q�҃���^��]á����   �AT�U�R�Ћu��P����a�������   �
�E�P�у���^��]�������������U����H��  ]��������������U����H��\  ]��������������U����H�U��t  ��V�uVR�E�P�у����S@���M��?����^��]�����U����H�U���  ��VWR�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]����������������U����H�U���  ��VWR�E�P�ы��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]����������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H�U�E��VWj R�UP�ERP��t  �U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�(_��^��]��U����H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    �����   j P�BV�Ћ����   �
�E�P�у�$��^��]���U����H��8  ]��������������U���  �\�3ŉE��M�EPQ������h   R连 ����|	=�  |#����H��0  hНhH  �҃��E� ���H��4  ������Rh��ЋM�3̓���  ��]�������U����H��  ��V�U�WR�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]����U����H��  ��V�U�WR�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]����U����H��p  ��$�҅�trh���M��)]�����P�E�R4Ph���M��ҡ��P�E�R4Ph���M���j �E�P�M�hicMCQ���������   ��M�Q�҃��M��]����]�U����H��p  ��$V�҅�u���H�u�QV�҃���^��]�Wh!���M��|\�����P�E�R4Ph!���M���j �E�P�M�hicMCQ���������   �QHP�ҋu�����H�QV�ҡ��H�QVW�ҡ����   ��U�R�Ѓ�$�M��=\��_��^��]������U����H��p  ��$V�҅�u���H�u�QV�҃���^��]�Wh����M��[�����P�E�R4Ph����M���j �E�P�M�hicMCQ���������   �QHP�ҋu�����H�QV�ҡ��H�QVW�ҡ����   ��U�R�Ѓ�$�M��m[��_��^��]������U����H��p  ��$�҅�u��]�Vh#���M���Z�����P�E�R4Ph#���M���j �E�P�M�hicMCQ����������   �Q8P�ҋ�����   ��U�R�Ѓ��M���Z����^��]���������������U����H��p  ��$�҅�u��]�Vhs���M��TZ�����P�E�R4Phs���M���j �E�P�M�hicMCQ�W��������   �Q8P�ҋ�����   ��U�R�Ѓ��M��5Z����^��]���������������U����H���  ]��������������U����H��@  ]��������������U����H���  ]��������������U��V�u���t���QP��D  �Ѓ��    ^]������U����H��H  ]��������������U����H��L  ]��������������U����H��P  ]��������������U����H��T  ]��������������U����H��X  ]��������������U����H��\  ]�������������̡��H��d  ��U����H��h  ]��������������U����H��l  ]�������������̡��H���  ��U����H�U���  ��VR�E�P�ыu��P���#X���M��;X����^��]�����U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H���  ]��������������U����H��l  ]��������������U����H���  ]��������������U����H���  ]��������������U����H��$  ]��������������U����H��(  ]��������������U����H��,  ]�������������̡��H��0  ����H��<  ��U����H���  ]�������������̡��H���  ��U����H���  ]������������������������������U����H��  ]�������������̡��H��P  ��U����H��`  ]�������������̡����   ���   ��Q��Y��������U����H�A�U��� R�Ћ��Q�Jj j��E�h�P�ыUR�E�P�M�Q��\�����B�P�M�Q�ҡ��H�A�U�R�Ћ��Q�J�E�P�у�,��]��h�PhD � �  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h�jhD �,�  ����t
�@��t]��3�]��������Vh�j\hD ����  ����t�@\��tV�Ѓ���^�����Vh�j`hD ����  ����t�@`��tV�Ѓ�^�������U��Vh�jdhD ���  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�jhhD ���Y  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh�jlhD ���  ����t�@l��tV�Ѓ�^�������U��Vh�h�   hD ����~  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h�   hD ���~  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�jphD ���I~  ����t�@p��t�MQV�Ѓ�^]� ��^]� ��U��Vh�jxhD ���	~  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�j|hD ����}  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�j|hD ���}  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� �������������U���Vh�h�   hD ���3}  ����t=���   ��t3�MQ�U�VR��h�j`hD �}  ����t�@`��t	�M�Q�Ѓ���^��]� �����̋���������������h�jhD �|  ����t	�@��t��3��������������U��V�u�> t+h�jhD �|  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h�jhD �A|  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�jhD ����{  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�jhD ���{  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�j hD ���|{  ����t�@ ��tV�Ѓ�^�3�^���Vh�j$hD ���L{  ����t�@$��tV�Ѓ�^�3�^���U��Vh�j(hD ���{  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�j,hD ����z  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�j(hD ���z  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�j4hD ���<z  ����t�@4��tV�Ѓ�^�3�^���U��Vh�j8hD ���	z  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�j<hD ���y  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh�jDhD ���|y  ����t�@D��tV�Ѓ�^�3�^���U��Vh�jHhD ���Iy  ����t�M�PHQV�҃�^]� U��Vh�jLhD ���y  ����u^]� �M�PLQV�҃�^]� �����������U��Vh�jPhD ����x  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�jThD ���x  ����u^Ë@TV�Ѓ�^���������U��Vh�jXhD ���ix  ����t�M�PXQV�҃�^]� U��Vh�h�   hD ���6x  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�h�   hD ����w  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�h�   hD ���w  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ���Vw  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ���w  ����u^]� �M���   QV�҃�^]� �����U��Vh�h�   hD ����v  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh�h�   hD �v  ����u���H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ��Q�u���BV�Ћ��Q�BVW�Ћ��Q�J�E�P�у�_��^��]��U��Vh�h�   hD ���v  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�h�   hD ���u  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   hD ���vu  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�h�   hD ���6u  ����t���   ��t�MQ����^]� 3�^]� �Vh�h�   hD ����t  ����t���   ��t��^��3�^����������������U��Vh�h�   hD ���t  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�h�   hD ���ft  ����t���   ��t�MQ����^]� ��������U��Vh�h�   hD ���&t  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh�h�   hD ����s  ����t���   ��t��^��3�^����������������VW��3����$    �h�jphD �s  ����t�@p��t	VW�Ѓ�����8 tF��_��^�������U��SW��3�V��    h�jphD �?s  ����t�@p��t	WS�Ѓ�����8 tqh�jphD �s  ����t�@p��t�MWQ�Ѓ������h�jphD ��r  ����t�@p��t	WS�Ѓ����V���������tG�]����E^��t�8��~=h�jphD �r  ����t�@p��t	WS�Ѓ�����8 u_�   []� _3�[]� ����������U��Vh�j\hD ���9r  ����t3�@\��t,V��h�jxhD �r  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�j\hD ����q  ����t3�@\��t,V��h�jdhD �q  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�j\hD ���vq  ����tG�@\��t@V�ЋEh�jdhD �E��E�    �E�    �@q  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�j\hD ����p  ����t\�@\��tUV��h�jdhD ��p  ����t�@d��t
�MQV�Ѓ�h�jhhD �p  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�j\hD ���ip  ������   �@\��t~V��h�jdhD �Cp  ����t�@d��t
�MQV�Ѓ�h�jhhD �p  ����t�@h��t
�URV�Ѓ�h�jhhD ��o  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh�jthD ���o  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�j`hD �~o  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh����_�����^��]� ������U���Vh�h�   hD �%o  ����tU���   ��tK�M�UQR�M�Q�Ћu��P������h�j`hD ��n  ����t%�@`��t�U�R�Ѓ���^��]ËE�uP���k�����^��]�����U���Vh�h�   hD ���n  ����tR���   ��tH�MQ�U�R���ЋuP������h�j`hD �Zn  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    �'�����^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t�����   P�B@��]� �E��t�����   P�BD��]� �����   R�PD��]� �����U����P@�Rd]�����������������U����P@�Rh]�����������������U����P@�Rl]�����������������U����P@�Rp]�����������������U������   ���   ]�����������U������   ���   ]����������̡��P@�Bt����̡��P@�Bx�����U����P@�R|]����������������̡��P@���   ������   �Bt��U����P@���   ]�������������̡��P@���   ��U����P@���   ]��������������U����P@���   ]��������������U����P@���   ]��������������U����P@���   ]��������������U����P@���   ]��������������U����P@���   ]��������������U���V��H@�QV�ҋM����t��#������Q@P�BV�Ѓ�^]� �̡��PH���   Q�Ѓ�������������U����P@�EPQ�JL�у�]� ���̡��P@�BHQ�Ѓ����������������U����P@�EP�EP�EPQ�J�у�]� ������������U����P@�EPQ�J�у�]� ����U����P@�EP�EPQ�J�у�]� U����P@�EPQ�J �у�]� ����U������   �R]��������������U������   �R]��������������U������   �R ]��������������U������   ���   ]�����������U������   ��D  ]�����������U����E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U������   ���   ]����������̡����   �B$����H@�Q0�����U����H@�A4j�URj �Ѓ�]����U����H@�A4j�URh   @�Ѓ�]�U����H@�U�E�I4RPj �у�]�̡��H|�������U��V�u���t���Q|P�B�Ѓ��    ^]��������̡��H|�Q �����U��V�u���t���Q|P�B(�Ѓ��    ^]��������̡��H@�Q0�����U��V�u���t���Q@P�B�Ѓ��    ^]���������U����H@���   ]��������������U��V�u���t���Q@P�B�Ѓ��    ^]��������̡��PH���   Q�Ѓ�������������U����PH�EPQ��d  �у�]� �U����H �IH]�����������������U��}qF uHV�u��t?�����   �BDW�}W���Ћ��Q@�B,W�Ћ��Q�M�Rp��VQ����_^]����������̡��P@�BT�����U����P@�RX]�����������������U����P@�R\]����������������̡��P@�B`�����U����H��T  ]��������������U����H@�U�A,SVWR�Ћ��Q@�J,���EP�ы��Z��h��hE  �΋��v;��Ph��hE  ���d;��P��T  �Ѓ�_^[]����U����PT�EP�EPQ�J�у�]� U����PT�EPQ�J�у�]� ����U����PT�EPQ�J�у�]� ����U����PT�E�R<��PQ�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U����HT�]��U����H@�AV�u�R�Ѓ��    ^]�������������̡��HT�hG  �҃�������������U����H@�AV�u�R�Ѓ��    ^]�������������̡��PD�BQ�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�BQ�Ѓ����������������U����PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U����PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U����PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U����PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U����PX�EPQ�J�у�]� ����U����PX�EPQ�J�у�]� ����U����PX�EPQ�J�у�]� ����U����PX�EPQ�J�у�]� ����U����PX�EPQ�J$�у�]� ����U����PX�EPQ�J �у�]� ����U����PD�EP�EPQ�J�у�]� U����HD�U�j R�Ѓ�]�������U����H@�AV�u�R�Ѓ��    ^]��������������U����HD�	]��U����H@�AV�u�R�Ѓ��    ^]��������������U����HD�U�j R�Ѓ�]�������U����H@�AV�u�R�Ѓ��    ^]��������������U����U�HD�Rh2  �Ѓ�]����U����H@�AV�u�R�Ѓ��    ^]��������������U����U�HD�RhO  �Ѓ�]����U����H@�AV�u�R�Ѓ��    ^]��������������U����U�HD�Rh'  �Ѓ�]����U����H@�AV�u�R�Ѓ��    ^]�������������̡��HD�j h�  �҃�����������U����H@�AV�u�R�Ѓ��    ^]�������������̡��HD�j h:  �҃�����������U����H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E������   �R�E�Pj�����#E���]�̡��HD�j h�F �҃�����������U����H@�AV�u�R�Ѓ��    ^]�������������̡��HD�j h�_ �҃�����������U����H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E����E�    ���   �R�E�Pj������؋�]� ̡��PD�B$Q�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ���������������̡��PD�B(Q�Ѓ���������������̡��PD�BQ�Ѓ����������������U����H �Ah]�����������������U����H@�AV�u�R�Ѓ��    ^]�������������̡��H �������U��V�u���t���Q P�B�Ѓ��    ^]���������U����P �EPQ�J4�у�]� ����U����P �EPQ�J�у�]� ����U����P �EPQ�J�у�]� ���̡��P �BQ��Y�U��V�uW�����//�����H �QVW�҃�_��^]� �����U����P �EPQ�J �у�]� ���̡��P �B,Q�Ѓ���������������̡��P �B0Q�Ѓ���������������̡��H\�������U����H\�AV�u�R�Ѓ��    ^]�������������̡��P\�BQ�Ѓ���������������̡��P\�BQ�Ѓ����������������U����P\�EPQ�J�у�]� ����U����P\�EP�EPQ�J�у�]� U����P\�EPQ�J�у�]� ���̡��P\�BQ�Ѓ����������������U����P\�EPQ�J �у�]� ����U����P\�EP�EPQ�J$�у�]� U����P\�EP�EP�EP�EPQ�J`�у�]� ��������U����P\�EPQ�J0�у�]� ����U����P\�EPQ�J@�у�]� ����U����P\�EPQ�JD�у�]� ����U����P\�EPQ�JH�у�]� ���̡��P\�B4Q�Ѓ����������������U����P\�EP�EPQ�J8�у�]� U����P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu���$�����H\�QV�҃���S���$��3���~B��I ���H\�U�R�U��EP�A`h���VR�ЋM��Q���$���U�R���x$��F;�|�_^[��]� ����������U���VW�}�E��P��� ���}� ��   ���Q\�BV�Ѓ��M�Q��� ���E���t]S3ۅ�~H�I �UR���e ���E�P���Z ���E;E�!�����Q\P�BV�ЋE@��;E��E~�C;]�|�[_�   ^��]� _�   ^��]� U����E�PH�B���$Q�Ѓ�]� ���������������U����PH�EPQ���   �у�]� �U����PH�EPQ���  �у�]� �U����PH�EPQ���  �у�]� �U����PH�EP�EPQ��  �у�]� �������������U����PH�EP�EPQ��  �у�]� ������������̡��PH���  Q�Ѓ�������������U����PH�EPQ���  �у�]� ̡��PH���   j Q�Ѓ�����������U����PH�EPj Q���   �у�]� ��������������̡��PH���   jQ�Ѓ�����������U����PH�EPjQ���   �у�]� ��������������̡��PH���   jQ�Ѓ����������U����PH�EPjQ���   �у�]� ���������������U����PH�EP�EPQ���   �у�]� �������������U����PH�EP�EPQ���   �у�]� ������������̡��PH���   Q�Ѓ�������������U����PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP��� ���������t�E���QH���   PVW�у���_^]� �����U��EVW���MPQ�,���������t�M���BH���   QVW�҃���_^]� ̡��PH���   Q�Ѓ������������̡��PH���   Q�Ѓ�������������U����PH�EPQ���   �у�]� �U����PH�EPQ���   �у�]� �U����PH�EP�EPQ��8  �у�]� �������������U����PH�EP�EPQ��   �у�]� ������������̡��PH���  Q�Ѓ������������̡��PH���  Q�Ѓ������������̡��PH���  Q�Ѓ������������̡��PH��  Q�Ѓ������������̡��PH��  Q�Ѓ�������������U����PH�EP�EPQ��  �у�]� �������������U����PH�EP�EP�EPQ��   �у�]� ���������U����PH�EP�EP�EP�EPQ��|  �у�]� �����U����PH�EPQ��  �у�]� ̡��PH��T  Q�Ѓ�������������U����PH�EP�EPQ��  �у�]� �������������U����PH�EPQ��8  �у�]� �U����PH�EPQ��<  �у�]� �U����PH�EP�EP�EPQ��@  �у�]� ���������U����PH�EPQ���  �у�]� ̡��PH��L  Q��Y��������������U����PH�EPQ��H  �у�]� ̡�V��H@�Q,WV�ҋ��Q��j �ȋ��   h�  �Ћ��QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡��P@�B,Q�Ћ��Q��j �ȋ��   h�  �������U����E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U����E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U����PH�EP�EP�EPQ��   �у�]� ��������̡��HH��  ��U����HH��  ]��������������U����E�PH��$  ���$Q�Ѓ�]� �����������̡��PH��(  Q�Ѓ�������������U����PH�EP�EPQ��,  �у�]� �������������U����E�PH�EP�E���$PQ��0  �у�]� ���̡��PH���  Q�Ѓ������������̡��PH��4  Q�Ѓ������������̋��     �������̡��PH���|  jP�у���������U����UV��HH��x  R��3Ƀ������^��]� ��̡��PH���|  j P�у��������̡��PH��P  Q�Ѓ������������̡��PH��T  Q�Ѓ������������̡��PH��X  Q�Ѓ�������������U����PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡��PH��`  Q�Ѓ�������������U����PH�EPQ��d  �у�]� �U����E�PH��h  ���$Q�Ѓ�]� ������������U����E�PH��t  ���$Q�Ѓ�]� ������������U����E�PH��l  ���$Q�Ѓ�]� ������������U����PH�EPQ��p  �у�]� �U����PH�EP�EP�EP�EPQ���  �у�]� �����U����PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U����E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E���HH�E���   R�U���$P�ERP�у�]����������������U���E�M� ��|�  �M;�|�M;�~��]�����������U����PH�E���   Q�MPQ�҃�]� ������������̡��PH���   Q��Y�������������̡��PH���   Q�Ѓ������������̡��PH���   Q��Y��������������U����PH�EP�EPQ���   �у�]� �������������U����PH�EP�EP�EP�EP�EPQ���  �у�]� ̡��PH��t  Q��Y�������������̋�� ,��@    ��,����Pl�A�JP��Y��������U���V��Hl�V�AR�ЋE����u
�   ^]� ���Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË��QlP�B�Ѓ�������U����Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E���HH�ER�U���$P���  R�Ѓ�]����U����HH���  ]��������������U����HH���  ]��������������U��U0�E(���HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U����HH���  ]��������������U����E�PH�EP���$Q���  �у�]� ��������U���V��������E����  �} ��   ���HH��p  SWj h�  V�ҋء��HH���   h�  V�]��ҋ������}����   �M3��u���������   �]�E�P�M�Q�MWV�z�����t^�u�;u�V������u�E�������L�;Ht-���Bl�S�@����QR�ЋD������t	�M�P�a���F;u�~��}�u�MF�u��)���;��u����E�_[^��]� 3�^��]� ������������U�����SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u���HH���  �'��u���HH���  ���uš��HH���  S�ҋȃ��E��t�W��������HH���   h�  S3��҃����  ���_�u����    ���Hl�U�B�IWP�ы�������   ���F�J\�UP�A,R�Ѓ���t�K�Q�M�������F�J\�UP�A,R�Ѓ���t�K�Q�M������E��;Pt&�F���Q\�J,P�EP�у���t	�MS�������v�B\�M�P,VQ�҃���t�M�CP�������QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U����HH���   ]�������������̡��PH���   Q��Y��������������U����HH���  ]��������������U�����P���   V�uW�}���$V�����E������At���E������z����؋��Q�B,���$V����_^]����������������U���0����U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١��]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U����HH�]��U����H@�AV�u�R�Ѓ��    ^]�������������̡��HH�h�  �҃�������������U����H@�AV�u�R�Ѓ��    ^]��������������U����HH�Vh  �ҋ�������   �EPh�  �P�������t]���QHj P���   V�ЋMQh(  �&�������t3���JH���   j PV�ҡ����   �B��j j���Ћ�^]á��H@�QV�҃�3�^]�������U����H@�AV�u�R�Ѓ��    ^]��������������U����HH�Vh�  �ҋ�����u^]á��HH�U�E��  RPV�у���u���B@�HV�у�3���^]�������U����H@�AV�u�R�Ѓ��    ^]��������������U����HH�I]�����������������U����H@�AV�u�R�Ѓ��    ^]��������������U����PH�EPQ���  �у�]� �U����PH�EPQ���  �у�]� ̡��PH���  Q�Ѓ�������������U����HH���  ]��������������U����E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡��PH���  Q�Ѓ�������������U����PH�EP�EPQ���  �у�]� ������������̡��PH��  Q�Ѓ�������������U����PH�EP�EP�EPQ���  �у�]� ��������̡��PH���  Q�Ѓ������������̡��PH���  Q�Ѓ�������������U����PH�EPQ��  �у�]� �U����PH�EPQ��  �у�]� ̋������������������������������̡��HH���  ��U����HH���  ]��������������U����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U����PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡��PH��,  Q�Ѓ�������������U����PH�EPQ��X  �у�]� ̡��PH��\  Q�Ѓ�������������U����HH��0  ]��������������U�����W���HH���   j h�  W�҃��} u�   _��]� Vh�  �������������   ���HH���   j VW�҃��M��������P�E�R0Ph�  �M����E���P�B,���$h�  �M��Ћ��Q@�J(j �E�PV�у��M�����^�   _��]� ^3�_��]� �����U��S�]�; VW��u7���U�HH���   RW�Ѓ���u���QH���   jW�Ѓ���t�   �����   ���QH���   W�Ѓ��} u(���E�QH�M���  P�ESQ�MPQW�҃��B�u��t;���U�HH�ER�USP���  VRW�Ћ����   �B(�����Ћ���uŃ; u���QH���   W�Ѓ���t3���   �W��u1���QH���   �Ћ��E�QH���   PW�у�_^[]� ���BH���   �у��} u0���M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ���QH�h  �Ћ؃���u_^[]� �����   �u�Bx���Ћ����   P�B|���Ѕ�tU���E�QH�MP�Ej Q���  VPW�у���t�����   �ȋBHS�Ћ����   �B(���Ћ���u�_^��[]� ��������������U��EV���u���HH���  �'��u���HH���  ���u���HH���  V�҃���u3�^]� P�EP���.���^]� ���������U���D���HH���   S�]VWh�  S�ҋ���HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��.
  �����   �B���Ћ�=�  ��  �QH���   Wh:  S�Ћ��QH�E����   h�  S�Ћ��QHW�����   h�  S�uԉ}��Ћ��QH�E苂  S�Ћ��QH�EЋ��  S�Ѓ�(�E��E�8���~~�M���M�I �MЅ�tMj�W�O  ���t@�@�Ẽ|� �4�~����%�������;�u/����Y  ;E�~�E؋��Y  E���E�;Pu�E���E��E�G;}�|��}� tv�u�j S�����������  ��������tV���a����}�;�uK���H���  �4�h@���h�  V�҃��E���N  �M�PVP�m���P�  ����}ܡ��H���  �4�h@���h�  V�҃��E����  �M�3�;�t;�tVQP��  ���E�;�~-���Qh@���h�  P���   �Ѓ��E�;���  ���E��QH��  j�PS�у�����  �u�;�tjS���������{  �������E���}���BH���   Wh�  S�у�3�9}ԉE�}��`  �}���}Ȑ�MЅ��R  �U�j�R�M  ����>  �M̍@�|� ���]�~����%�������9E���  ���W  �E�3�3�9C�E܉M���   ��$    �����������tk�]��}������������ϋ9�<��}�@�҉��y�]��|��]�@@�z�<��y�]��|��]�@@�z�<��I�}��]�@���M��}�@����@�M�A;K�M��t����E؅��9  �+U�j��PR�M��:  �M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$���U����4�"�M����t��U����t�
�M����t�M���;]�|��E܃�F;]؉M��	����U�;U��
  �U�R��o���E�P�o���M�Q�o����_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���P�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@��;EԉE��}�������U�R�m���E�P�m�����  ���   �B����=  ��  ���QH���   j h(  S�Ћ��QH�����   h(  S�ЋЃ�3��U؅�~'����    �ǅ�t�|� t�4N��tN�@;�|�u��u܋��Q���  �4v�h@���hK  V�Ѓ��E�����   �M��t��tVQP���  ���u؋��Q���  �h@���hP  V�Ѓ��E���tP��t��tVWP趤  ���M����+��RH��PQ�E���   S�Ѓ���u�M�Q�Rl���U�R�Il����_^3�[��]á��HH���   j h�  S�҉E����HH���   j h(  S��3�3���3�9]؉E��}ĉ]��7  �U��څ��  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�F@F����;�|��}ă|� ts�U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�F�v�Ћ��A�B�A�B�A�B�A�B�I�J�U�F<ډ}�C;]؉]�������M�3�3�;�~�U����$    ��t���   @;�|��U�R�j�����E�P�{j����_^�   [��]�/�:�F�R�������������U��U��t�M��t�E��tPRQ�`�  ��]������������U��E� �M+]� ���������������U��V��V�,����Hl�AR�Ѓ��Et	V�m������^]� ����������h�Ph�f �.  ���������������U���Vh�h�   h�f ���S.  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh�h�   h�f ����-  ����t���   ��t�M�UQ�MRQ����^]� U���Vh�h�   h�f ���-  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh�h�   h�f ����,  ����t���   ��t�M�UQ�MRQ����^]� U��Qh�h�   h�f �,  ����t���   �E���t�EP�U�����]��P���]�������������U���h�h�   h�f �f,  3Ƀ�;�tK9��   tC�E���   ���M��$Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]ËE�   � �  �P�P�H�H�H��]��U��h�h�   h�f ��+  ����t���   ��t]��]����U��h�h�   h�f �+  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h�h�   h�f �I+  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h�h�   h�f ��*  ����t���   ��t]��3�]��U���Vh�h�   h�f �*  ����tZ���   ��tP�M�UWQR�M�Q�Ћ��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]á��H�u�QV�҃���^��]����������h�h�   h�f �*  ����t���   ��t��3��������U��h�h�   h�f ��)  ����t���   ��t]��]����U��VWh�h�   h�f �)  ������tb���    tY�E �M�UP��Q�HR�Q����V�ҡ��H�A�UVR�Ћ��   ���ы����B�P�MQ�҃� ��_^]á��H�A�UR�Ѓ�_3�^]���U��VWh�h�   h�f �)  ������tb���    tY�E �M�UP��Q�HR�Q����V�ҡ��H�A�UVR�Ћ��   ���ы����B�P�MQ�҃� ��_^]á��H�A�UR�Ѓ�_3�^]���U���Vh�h�   h�f �u(  ����tZ���   ��tP�M�UWQR�M�Q�Ћ��u���B�HV�ы��B�HVW�ы��B�P�M�Q�҃�_��^��]á��H�u�QV�҃���^��]����������U���Vh�h�   h�f ��'  ����tS���   ��tI�MWQ�U�R�Ћu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]Ë��Q�u�BV�Ѓ���^��]����������������U���Vh�h�   h�f �5'  ����tS���   ��tI�MWQ�U�R�Ћu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]Ë��Q�u�BV�Ѓ���^��]����������������U��h�h�   h�f �&  ����t���   ��t]��]����U��h�h�   h�f �i&  ����t���   ��t]��]����U��M��U+u&�A+Bu�A+Bu�A+Bu�A+Bu�A+B]����������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���h��   h�   h�f �E��  �E��E��E�    �E�    �E�    ��#  ����t���   ��t	�M�Q�Ѓ��UR�E�P��������]��U��E��u���MP�EPQ�c�����]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h��j;hj�b������t
W���^����3��F��u_^]� �~ t3�9_��^]� ���H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ���H<�Q��3Ʌ����^��������������̃y t�   ËA��uË��R<P��JP�у��������U����u���H�]� ���J<�URP�A�Ѓ�]� ���������������U�����u���H�]Ë��J<�URP�A�Ѓ�]�U�����$V��u���H�1����J<�URP�A�Ѓ������Q�J�E�SP�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h̞P�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���[t.���B�u�HV�ы��B�P�M�Q�҃���^��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�u�QV�ҡ��H�A�U�VR�Ћ��Q�J�E�P�у���^��]���������������U�����$SV��u���H�1����J<�URP�A�Ѓ������Q�J�E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h̞P�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���t/���B�u�HV�ы��B�P�M�Q�҃���^[��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h̞P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у����3������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�u�QV�ҡ��H�A�U�VR�Ћ��Q�J�E�P�у���^[��]����������������U�����$SV��u���H�1����J<�URP�A�Ѓ������Q�J�E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h̞P�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���t/���B�u�HV�ы��B�P�M�Q�҃���^[��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h̞P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у����3������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h̞P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у�����������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҋu�E�P���#p�����Q�J�E�P�у���^[��]�������U�����$SV��u���H�1����J<�URP�A�Ѓ������Q�J�E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Jj j��E�h̞P�ы��B�@@�� j �M�Q�U�R�M��Ћ��Q�J���E�P���у���t/���B�u�HV�ы��B�P�M�Q�҃���^[��]á��P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h̞P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у����3������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M��ҡ��H�A�U�R�Ћ��Q�Jj j��E�h̞P�ы��B�@@��j �M�Q�U�R�M��Ћ��Q�J���E�P���у�����������P�E��RHjP�M��ҡ��P�E�M��RLj�j�PQ�M���j h̞�M���m�����P�R@j �E�P�M�Q�M��҅����H�A�U�R���Ѓ���t/���Q�u�BV�Ћ��Q�J�E�P�у���^[��]Ë��M��B�PHjQ�M��ҡ��P�E�M��RLj�j�PQ�M��ҋu�E�P����l�����Q�J�E�P�у���^[��]���������������U����H<�A]����������������̡��H<�Q�����V��~ u>���t���Q<P�B�Ѓ��    W�~��t�������W��V�����F    _^��������U���V�E�P���������P��������M��������^��]��̃=� uK����t���Q<P�B�Ѓ���    ����tV���@���V�ZV������    ^������������U���8���H�AS�U�V3�R�]��Ћ��Q�JSj��E�hОP�ы��B<�P�M�Q�ҋ���H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��  �M�Q�U�R�M���  ����   W�}�}���   �����   �U��ATR�Ћ�����tB���Q�J�E�P���у��U�Rj�E�P���<k�����Q�ȋBxW���E���t�E� ��t���Q�J�E�P����у���t���B�P�M�Q����҃��}� u"�E�P�M�Q�M��/  ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3ۉ]�;�u_���H�A�U�R�Ћ��Q�JSj��E�hОP�ы��B<�P�M�Q�ҋ���H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��!  �M�Q�U�R�M��q  ���p  W�}��I �E����   �����   �U��ATR�Ћ�������   ���Q�J�E�P���ы��B���   ���M�Qj�U�R���Ћ��Q�J���E�P�ы��B�P�M�QV�ҡ��H�A�U�R�Ћ��Q�Bx��W�M����E��t�E ��t���Q�J�E�P����у���t���B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*�����   P�BH�Ћ��Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��s  �EP�M�Q�M�u��u�  ����   �u���E���tA��t<��uZ�����   �M�PHQ�ҋ��Q���ȋBxV�Ѕ�u-�   ^��]Ë����   �E�JTP��VP�[�������uӍUR�E�P�M��4  ��u�3�^��]����������V��~ u>���t���Q<P�B�Ѓ��    W�~��t������W�Q�����F    _^�������̋�� ����������������������̅�t��j�����̡��P��  ����P��(  ��U����P��   ��V�E�P�ҋuP�������M��������^��]� ��������̡��P��$  ��U����H��  ]��������������U����H���  ]�������������̡��H��  ��U����H���  ]��������������U����H��x  ]��������������U����H��|  ]�������������̡��H��d  ��U����H��p  ]��������������U����H��t  ]��������������U���EV�����t	V��O������^]� �������������̸   � �������̸   @� �������̸   � �������̸   � ��������U����H�QV�uV�҃���^]� �3�� �����������3�� �����������3�� �����������U����   h�   ��@���j P�$d  �M�Eh�   ��@���R�M��MPQjǅ`���    �9x���� ��]���U����   V�u��u3�^��]�h�   ��@���j P��c  �M�U�Eh�   �M���@���Q�U��U��@����ERPj��`���ǅD��� ��E�б�E� ��E� ��E�0��E�P��E���E���E�@��w���� ^��]������U���   SV�u(3ۉ]���u���H�A�UR�Ѓ�^3�[��]Ë��Q�B<W�M3��Ѕ��'  �l8  �E���tq�MQ�M��)���Wh��M��[c��P�M������u�Wj��U�R�E�P��\���Q�_?�������P��x���R�������P�E�P������P���9  �E���t�E� �� t�M�����0�����t��x������������t��\�������
�����t�M̃���������t���Q�J�E�P����у���t�M�������}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R�_7  ����E$�M�UVP�Ej QRP������������Q�J�EP�у���_^[��]���������������̋�`����������̋�` ����������̋�`����������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V���5  �����   �ESP�M��x������Q�J�E�P�ы��B�Pj j��M�h�Q�҃��E�P�M��<���j j��M�Q�U�R��d���P������P�M�Q�������P�U�R��������P��6  ���M����q����M��i�����d����^����M��V������H�A�U�R�Ѓ��M��:�����[t	V��4  ����^��]� ���U��EVP���?  �����^]� �����Q�4  Y���������U��E�M�U�H4�M�P �U��M�@ ��@8б�@<��@@@��@D ��@H ��@L��@P0��@l��@X`��@\���@`@��@d ��@TP��@h0��@p���@t���P0�H(�@,    ]��������������U���   h�   ��`���j P�T^  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�Ur����8��]��������������̋�`<����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`,�����������U��E��u�E�M���   ]� �����������U��EHV����   �$����   ^]á@���uT�EP�g�����=�2  }�����^]Ëu��t�h�jmhj�KH������t ���m���� ��tV���|����   ^]��     �   ^]ËM�UQR�5����������H^]�^]�����-u.�����}���� ��t������V�G�����     �   ^]Ã��^]ÍI ��Y�`�����>�U���EV���V��������Au���H��0  h0�j,�����^��^]� �����U���W������G���U�� �������A�  ������A��   ���������AuR������AuKV���[y  ���Ty  �ȅ�u��^����__��]Ëƙ����ʅ�u�u��E�^������__��]���������Au������=x���������Au6�����������U������G�����_��������Au�����U����_�
����������=  �E����U������������A{���������__��]�������������__��]����U�����V�E��������At�����������Au��������������$��v  ���������^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3������;���W���$���v  ��E������$�lv  �V����������Au���H��0  h0�j�����^����_u������������^]� ���U������EV�ы�������z!���؋H��0  h0�j5�����U������$��u  �]��F�$��u  �}��$��u  ��E�$�u  �^�����&���^��]� ���������������U������   �BXQ�Ѓ���u]� ���Q|�M�RQ�MQP�҃�]� ���U������   �BXQ�Ѓ���u]� ���Q|�M�R8Q�MQP�҃�]� ���U��EV��j ����Qj j P�B�ЉF����^]� ��̡�Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ���Q�MP�EP�Q�JP�у��F�   ^]� ����U��M��P]����U��M��P]����U��M��P]����V������F    ���HP�h0�Vh �h��҉F����^����������̃y ���u���PP�A�JP��Y��U��A��u]� ���QP�M�Rj Q�MQP�҃�]� ��U��A��t���QP�M�RQP�҃�]� ������������U��A��t���QP�M�RQP�҃�]� �����������̡��HP���   ��U����HP���   ]�������������̡��HP�QP�����U����HP�AT]����������������̋��     �@    �V����t)���QPP�BL�Ћ��QP��J<P�у��    ^�������������U��SV�ً3�W;�t���QPP�B<�Ѓ��3�s�}�Eh0�W�C���QP�J8h �h�P�EP�у�9u�~M�I ���z u!���@   ���QP���H�RQ�҃����HP��A@VR�Ћ�F��;u�A|�3�9_^��[]� ��������U��SVW��3�9w~<�]���HP��A@VR�Ѓ���t-���QPj SjP�B�Ѓ���tF;w|�_^�   []� ���QP��JLP�у�_^3�[]� �����������̡��PP��JDP�у�������������̡��PP��JHP��Y��������������̡��PP��JLP��Y���������������U��U�E�@R�URP�I���]� �����U��V��~ ���u���HP�V�AR�Ѓ��Et	V�>������^]� ����U��E�M�UP��P�EjP�l����]��������������̸   �����������U��V�u��t���u6�EjP�l������u3�^]Ë��m����t���t��U3�;P��I#�^]�������U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �������������U��V�u�F��F�����������������\q  ����������D�Ez��^��P�X]��������������N�X�N^�X]��������P�P�P�P �P(�P0�P8�P@�PH�PP�PX����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��5�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A �A�A(�A�������������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E������X�X]� ̋�3ɉ�H�H�H�V��V�W0���FP�N0��3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  S�]���q  ��؋�U��M�U�>�U��@�����@�U��@�B�@�������@���@�   ;����U��p  �w�����  �w�������F�B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]؋�R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ɍU��R�[�[������E��KH��P�E�SL��H�щKP�P�ST�H�KX�P�����S\��z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����M��}������3�3����u��u�|+�A�����B�4�u�0u��u�p�����u�u�U�E;�}�Q���E����U��U��1���@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���@�D��KX�@�U�����]��C���@�K0���@�KH���C ��C�@�K8���@�KP���C(��C�C@�H���@3����KX���U��r  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������]��E�E����]���E����]��E׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���@�   �KXE)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� ������������hPh_� �������������������hjh_� ��������uË@����U��V�u�> t/hjh_� �c�������t��U�M�@R�Ѓ��    ^]���U��Vhjh_� ���)�������t�@��t�MQ����^]� 3�^]� �������U��Vhjh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vhjh_� ����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vhjh_� ���Y�������t�@��t�MQ����^]� 3�^]� �������U��Vhj h_� ����������t�@ ��t�MQ����^]� 3�^]� �������U��Vhj$h_� �����������t�@$��t�MQ����^]� 2�^]� �������Vhj(h_� ����������t�@(��t��^��3�^������Vhj,h_� ���l�������t�@,��t��^��3�^������U��Vhj0h_� ���9�������t�@0��t�MQ����^]� 3�^]� �������U��Vhj4h_� �����������t�@4��t�M�UQR����^]� ���^]� ��Vhj8h_� ����������t�@8��t��^��3�^������U��Vhj<h_� ����������t�@<��t�MQ����^]� ��������������U��Vhj@h_� ���I�������t�@@��t�MQ����^]� ��������������U��VhjDh_� ���	�������t�@D��t�MQ����^]� 3�^]� �������U��VhjHh_� �����������t�@H��t�MQ����^]� ��������������VhjLh_� ����������t�@L��t��^��3�^������VhjPh_� ���\�������t�@P��t��^��3�^������VhjTh_� ���,�������t�@T��t��^��^��������VhjXh_� �����������t�@X��t��^��^��������Vhj\h_� �����������t�@\��t��^��^��������U��Vhj`h_� ����������t�@`��t�M�UQR����^]� 3�^]� ���U��Vhjdh_� ���Y�������t�@d��t�M�UQR����^]� 3�^]� ���U��Vhjhh_� ����������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vhjlh_� �����������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vhjph_� ���y�������t�@p��t�M�UQR����^]� 3�^]� ���U��Vhjth_� ���9�������t�@t��t�M�UQR����^]� 3�^]� ���U��Vhjxh_� �����������t�@x��t�M�UQR����^]� 3�^]� ���U��Vhj|h_� ����������t�@|��t�MQ����^]� 3�^]� �������U��Vhh�   h_� ���v�������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vhh�   h_� ���&�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vhh�   h_� �����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vhh�   h_� ���f�������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vhh�   h_� ����������t���   ��t�MQ����^]� 3�^]� �U��Vhh�   h_� �����������t���   ��t�MQ����^]� ��������U��Vhh�   h_� ����������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vhh�   h_� ���F�������t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E����������m������U�_��^�U�[���U������������������������Y  ����������D�Ez����P�X��]� �������E�����E����X�M��X��]� �����U���@����A���E�    �����]��]��]�����������]��]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P�q����F�@��R�M��_����~���Q�M��M����v;�t�v��P�M��7����M����m��M�u�_^[�M�UQR�M��������]� ��������������̋Q3���|�	��t��~�    t@����u��3���������U��QV�u;��}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��|+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~#V�1�d$ ���   @u	�����t@����u�^���̋QV3���~�	�d$ ����ШtF����u��^���������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%���;��E���}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$����E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ��b�x�����������U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�����FP����3����F�F^��U��SV��WV����^S����E3����~�~;�t_���Q���   h����jIP�у��;�t9�}��t;���B���   h����    jNQ�҃����uV�;����_^3�[]� �E�~_�F^�   []� ����������U��SV��WV����^S�����}3Ƀ��N�N;���   9��   �G;���   ���Q���  h����jlP�у����t=� t@�G��t9���Jh����    ���  jqR�Ѓ����u������_^3�[]� �O�N�G�Q��    R�F�QP����������t�N�WP��QPR�ث����_^�   []� ���������U��SV��WV����~W����3Ƀ��N�N9M��   �E;���   ��    ���H���  h��h�   S�҃����t=�} tH�E��tA���Q���  h����h�   P�у����u������_^3�[]� �U�V�,�F   ���H���  h��h�   j�҃����t��E�M�F�PSPQ�Ѫ���E����t!�V�?�W�RWP赪����_^�   []� ��M�_^�   []� ���U��Q�A�E� ��~LS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U�����u�_^[�E��Ћ�]� ���������U��S�]V��3�W�~���F�F�CV;C��   �D��W�>��3��F�F���Q���   h��jIj�Ѓ������   ���Q���   h��jNj�Ѓ����uV������_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� ���W���3��F�F���B���   h��jIj�у����t[���B���   h��jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP��������^]� ���������̡��H���   ��U����H���   V�u�R�Ѓ��    ^]����������̡��P���   Q�Ѓ�������������U����P�EPQ���   �у�]� ̡��H�������U����H�AV�u�R�Ѓ��    ^]��������������U����H�AV�u�R�Ѓ��    ^]��������������U����P��Vh�  Q���   �E�P�ы����   �Q8P�ҋ�����   ��U�R�Ѓ���^��]��������������̡��P�BQ�Ѓ����������������U����P�EPQ�J\�у�]� ����U����P�EP�EP�EP�EP�EPQ���   �у�]� �U����P�EP�EP�EP�EPQ�JX�у�]� �������̡��P�B Q��Y�U����P�EP�EP�EP�EPQ���   �у�]� �����U����P�EP�EP�EPQ�J�у�]� ������������U����H��   ]��������������U����P�R$]�����������������U����P��x  ]�������������̡��P��|  ��U����P�EP�EP�EP�EPQ�J(�у�]� ��������U����P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U����P�EP�EP�EP�EPQ�J,�у�]� ��������U���V��H�QWV�ҋ����H�QV�ҋ��Q�M�R4Q�MQ�MQOWHPj j V�҃�(_^]� ���������������U����P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U����P�EP�EPQ�J@�у�]� U����P�EPQ�JD�у�]� ���̡��P�BLQ�Ѓ���������������̡��P�BLQ�Ѓ���������������̡��P�BPQ�Ѓ����������������U����P�EPQ�JT�у�]� ����U����P�EPQ�JT�у�]� ����U����P�EP�EPQ���   �у�]� �������������U����P�E���   ��VP�EPQ�M�Q�ҋu�    �F    �����   j P�BV�Ћ����   �
�E�P�у� ��^��]� ������̡��P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡��H�������U����H�AV�u�R�Ѓ��    ^]��������������U����P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U����P�EPQ�J�у�]� ���̡��P�BQ��Y�U����P�EP�EPQ�J�у�]� U��VW��褽���M�U�x@�EPQR��莽���H ���_^]� �U��VW���t����M�U�xD�EPQR���^����H ���_^]� �V���H����xH u3�^�W���6����΍xH�,����H �_^�����U��V�������xL u3�^]� W��� ����M�U�xL�EPQR�������H ���_^]� �������������U��V���ż���xP u���^]� W��诼���M�U�xP�EP�EQRP��蕼���H ���_^]� ��������U��V���u����xT u���^]� W���_����M�xT�EPQ���M����H ���_^]� U��V���5����xX u���^]� W�������xX�EP�������H ���_^]� ����U���S�]VW���t.�M�覢�����߻���xL�E�P���ѻ���H ��ҍM������}��tZ���H�A�U�R�Ћ��Q�J�E�WP�ы��B�P�M�Q�҃����y����@@��t���QWP�B�Ѓ�_^[��]� ������U��V���E����x` u
� }  ^]� W���-����x`�EP�������H ���_^]� ��U��VW�������xH�EP��������H ���_^]� ���������U��SVW���Ӻ���x` u� }  �#��迺���x`�E���P��謺���H ��ҋ����H�]�QS�҃�;�A���H�QS�҃�;�,���o����M�U�xD�EPQSR���X����H ���_^[]� _^�����[]� ��������������U��V���%����xP u
�����^]� W�������M�U�xP�EP�EQ�MR�UPQR�������H ���_^]� ��������������U��V���Ź���xT u
�����^]� W��譹���M�xT�EPQ��蛹���H ���_^]� ��������������U��V���u����xX tW���g����xX�EP���Y����H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u���  ����t.�E�;�t'���J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡��H��   ��U����H��$  V�u�R�Ѓ��    ^]�����������U����UV��H��(  VR�Ѓ���^]� �����������U����P�EQ��,  P�у�]� �U����P�EQ��,  P�у����@]� �����������̡��H��0  ����H��4  ����H��p  ����H��t  ��U��E��t�@�3����RP��8  Q�Ѓ�]� �����U����P�EPQ��<  �у�]� �U����P�EP�EP�EPQ��@  �у�]� ���������U����P�EP�EPQ��D  �у�]� �������������U����P�EPQ��H  �у�]� �U����P�E��L  ��VWPQ�M�Q�ҋu�����H�QV�ҡ��H�QVW�ҡ��H�A�U�R�Ѓ�_��^��]� ��������������̡��P��T  Q�Ѓ�������������U����P�EPQ��l  �у�]� ̡��P��P  Q�Ѓ�������������U����P�EPQ��X  �у�]� ̡��H��\  ��U����H��`  V�u�R�Ѓ��    ^]�����������U����P�EP�EP�EP�EP�EPQ��d  �у�]� �U����P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w���y����3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7�������xP t$S������j j �XPj�FP���ʹ���H ���[�    �~` t���H�V`�AR�Ѓ��F`    _^������������U��SV��Fx���Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR�3������u#���h ����H��0  h  �҃��E�~P���l|���j j jW�����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ���Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ��i����F|��u�E�~x��t�    �F`_^]� �M�Fx������t�3�_^]� U��QVW�}����>  ���H�QhV�҃�����u"�H��0  h �h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���  �EF;u�|�UR�} ����_�   ^��]� �������������U��QVW�}����~  ���H�QhV�҃�����u"�H��0  h �h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'�����QP�Bh�Ѓ���t�M��R���,  F;u�|ʍEP������_�   ^��]� �������������h �h�   hh�   �g������t�������3��������V���(����N^�_v�����������������U��VW�}�7��t��������N�3v��V�M�����    _^]�hPh�f ��������������������U��hjh�f ��������t
�@��t]�����]�������U��Vhjh�f �k���������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�Ju���E�NP�у�4�M���tu����^]ÍM�gu�����^]��U��hjh�f ���������t
�@��t]��3�]��������U��hjh�f ���������t�x t�P]��3�]������V��FW��u�~��N�<��u�< ��u_3�^á��H�F��  hP�j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� }(�V;Vu��������t�F�N��    �F9~|؋V;Vu���������t��F�N�U���F_�   ^]� ��������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T����H;ǉ�F�M���F_�   ^]� ����U��E��|2�Q;�}+J;Q}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�����3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�A�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W��������3����_�F�F^��������������U���SV�uW���^S�}�����3���F�F�O�N�W���V9G�E~|��I �O���F�U�9FuL��u�~��~��t���< ��tY���H���  hP�j8��    RP�у���t0�~�}���V��M����E�F@;G�E|�_^�   [��]� _^3�[��]� U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|���P�����_^]� �U����E�Qj�E��ARP�M��E����+�����]� �����U����Q�Ej�E��A�MRPQ�M��E����G�����]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q�L���t!�A��t�B�A�Q�P�A    �A    �̋�� ���@L��HV3��q�q�P�r�r�L��p�p�p�P�H^������V����������F3��FL�;�t�N;�t�H�F�N�H�V�V�F�FL�;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3��L�;�t�F;�t�A�F�N�H�V�V�Et	V��������^]� ������������U��V��W�~W�������3����E��F�Ft	V�A�����_��^]� ������U��V��������Et	V��������^]� ��U���V�u��u��=  �@�E���=  ���E�F�}� �E�u�E�H�����   �� ��   S�]W�   ;�s��uS�7  Y��u�   �F�Xt}��u�]��}��7  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPW�u�j �c6  ��$��u������E�t	�M����_[^�Ë�U��V��<  �@�u��<  jh   �F�==  YY�F��th   �L6  P�v�,  ���F   ��26  �f �F��^]Ë�Wh8�������uV� V��  �����Y|�^��_�h8�����}V� V�  �����Y|�^Ë�U��E��V��}k� P�  Y��^]� ���}k� P�  YË�U���u�x0  Y��t]��=  ]ËI�������t�j���Ë�U��V��������EtV�����Y��^]� ��U��E���t趕����t�j���]Ë�U��Qj �M��@���h�������%� Y�M��N����á�Ë�U��=� uh�����  Y�E��]�j���C>  j �M�������}�e� �w��GN���8 t�������t�j�����w��w�b  �M��Y�M�������Y>  Ë�U��Qj �M�������ȋ j�����������u�M������Ë�U��=� uh�����Yj����Y��t����M�H�3���]Ë�U��E�xP v�xTr�@@���@Pj �L  YY]�j�6��H=  ��u��F   3��E��F�F�F�Eh���N����F�r �����w=  � j�d���<  ��u����V�E�   ����Yj j�N�7������8=  Ë�U��V�������EtV����Y��^]� j����<  ������u{P�M��2�����!u�����uXj4�e���Y�ȉM��E���t
V�������3�V�E� ������N�F?   �$���+���Ή5�����������M���M���������}<  Ë�U��E�xVWr�p��pj j �J  YY��u����}P�O<������tVj �J  YY��u���P�OX���_^]Ë�U��VW���w ��vW�u�V�6����u�_^]� ��U��V�uWj ��������F��t�8P�[���Y�ǅ�u�F �f ��t�8P�A���Y�ǅ�u�f  _^]Ë�U��V�u�~ v�F����F��� V����Y�N$��tj����^]Ë�Vj�������P��2  YY��^Ë�V���6�0  �6�����YY^��1�.  Y��1�5  YË�U���V�u��u�7  �@�E��d7  ���E�F�}� �E�u�E�H�����   �� ��   S�]��   s!��uS��1  Y��u�   �F�X��   ��u�]��}��0  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPh   �u�j �0  ��$��u������E�t	�M����[^�Ë�U��V�u������Ƞ��^]� �Ƞ�i����U��V���Ƞ�V���EtV�Z���Y��^]� jD����Y9  hР�M�����e� �E�P�M�����h(��E�P�B  �jD����!9  h��M��q���e� �E�P�M��P���hx��E�P�
  ̋�U��V�u���B#���Ƞ��^]� ��U��USVW�ڋ�����   ��@t����t��3Ɂ�;���3�A;�t�� �@��u��������� u3��^��t%��t �uh���u�H  ����t	P�  Y���u����V�u�wH  ������t���tjj V�8  ����tV�ŋ�_^[]Ë�U���  �\�3ŉE��Eh  Ph  ������Pj �K  ����t3���u�������uP��������M�3��  �Ë�U���u� �]Ë�U���u�$�]Ë�U���u�(�]Ë�U���u�,�]Ë�U������u]�76  �MH�����]����@�����t�������
r������̋L$WSV��|$��to�q��tU���L$���:�t��t���:�t
��u�^[_3�Ê��:�u�~��a��t(���:�u��A��t�f���:�t��3�^[_���J  �G�^[_Ë�^[_Ë�Q����:K  YË�U��V��������EtV�q���Y��^]� ��U��E��	Q��	P�tK  ��Y�Y@]� ��U��E��t���8��  uP�  Y]Ë�U��EV���F ��uc�cU  �F�Hl��Hh�N�;�t�0��Hpu�N9  ��F;8�t�F�0��Hpu�M  �F�F�@pu�Hp�F�
���@�F��^]� ��U����\�3ŉE�S3�V;�u�xX  j^SSSSS�0�e  ���5  �uW��W  YY;Er��ЋU��H;�u ��8t�<a|<z, �A8u�3���   j�p�   SSj�WVQR�T+  �ȃ�$�M�;�u��W  � *   ��W  � �   9Ms���W  j"�^���;�~Ej�3�X���r9�A=   w� X  ��;�t� ��  �P��   Y;�t	� ��  ���M�E���]�9]�u�~W  �    냋U�j�pQ�u�j�WV�pR�*  ��$��t�u��uW��   ������<W  j*Y����u������Y�ƍe�^[�M�3��  �Ë�U���W�u�M�������}�E�P�u�_����}� YY_t�M��ap��Ë�U��j �u�u������]Ë�U��S3�9duA�E;�u�V  SSSSS�    �	  ��3��/��8t)�
��a|
��z�� �
B8u��Sj��u�X����E��[]Ë�U��MS3�VW;�t�};�w�KV  j^�0SSSSS�8	  �����0�u;�u��ڋъ�BF:�tOu�;�u��V  j"Y�����3�_^[]�;\�u���hV  �����������̋T$�L$��ti3��D$��u��   r�=�+ t�W  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�ø_s������Fj����i���3j����i�������r����i���i����hË�U�������c  �} �@t�	c  ��]���U��WV�u�M�}�����;�v;���  ��   r�=�+ tWV����;�^_u^_]��c  ��   u������r*��$���Ǻ   ��r����$�(�$�$��$���8d�#ъ��F�G�F���G������r���$��I #ъ��F���G������r���$��#ъ���������r���$��I ��������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���$,8L�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�������$�`�I �Ǻ   ��r��+��$���$������F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I dlt|�����D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$���������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ���` �` � ��Ë�U��S�]VW��������t&P�l,  ��FV�-  YY�G��t�3VP��������g �G   ��_^[]� ��U��S�]V������C�F���CWt1��t'P�,  ��GW��  YY�F��t�sWP�/������	�f ��F_��^[]� �y ���t	�q��  YËA��u���Ë�U��V�EP�����������^]� ��U��V�u���R��������^]� ���������U��V�������EtV�	���Y��^]� ��U��V������c����EtV�����Y��^]� ��U��V�uW3�;�u3��e9}u�O  j^�0WWWWW�  �����E9}t9urV�u�u�  �����uW�u������9}t�9us�bO  j"Y����jX_^]�������������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[Ë�U��EVW3�;�tG9}u�~N  j^�0WWWWW�k  �����)9}t�9Es�YN  j"Y�����P�u�u�_�����3�_^]Ë�U��E�D]Ë�U���(  �\�3ŉE������� SjL������j P������������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������@�j ���<���(���P�8���u��uj�>]  Yh ��4�P�0��M�3�[�����Ë�U���5D�G  Y��t]��j��\  Y]����3�PPPPP�������Ë�U��� �EVWjY�ȡ�}��E��E_�E�^��t� t�E� @��E�P�u��u��u��D��� jh���i  �u��tu�=|+uCj�^  Y�e� V��^  Y�E��t	VP��^  YY�E������   �}� u7�u�
j�]  Y�Vj �5��L���u�L  ���H�P�K  �Y�ui  Ë�U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$����U��QQSVWd�5    �u��E��j �u�u��u�o �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�;v  �� �E�_^[�E���]Ë�U��V��u�N3�����j V�v�vj �u�v�u��u  �� ^]Ë�U���8S�}#  u�2�M�3�@�   �e� �E�^�\��M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E���F  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M�����E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u��t  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����-���u�u  �M�N��k���M9H};H~���u	�M�]�u�} }ʋEF�0�E�;_w;�v�Lu  ��k�E�_^[�Ë�U��EV�u��]E  ���   �F�OE  ���   ��^]Ë�U���:E  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V�E  �u;��   u�E  �N���   ^]���D  ���   �	�H;�t���x u�^]�t  �N�H�ҋ�U����\��e� �M�3��M�E��E�E�E@�E�T�M��E�d�    �E�E�d�    �uQ�u�t  �ȋE�d�    ����jh���=e  3��}�3��u;���;�u ��G  �    WWWWW�����������   V�gu  Y�}��F@uwV�z  Y���t���t�����ȃ����@����A$u)���t���t���������@����@$�t�_G  �    WWWWW�K������M��9}�u�Nx
��A��V�u  Y�E��E������   �E��d  ËuV�u  Y�jh���9d  3��}�3��u;���;�u ��F  �    WWWWW�����������   V�ct  Y�}��F@uwV��x  Y���t���t�����ȃ����@����A$u)���t���t���������@����@$�t�[F  �    WWWWW�G������M��9}�u!�Nx��E�����V�u�x  YY�E��E������   �E��c  ËuV�t  YË�U��V�u�F@WuyV�1x  Y�����t���t�ȃ��������@����A$u&���t���t�ȃ������@����@$�t�E  3�WWWWW�    �y���������JS�]���t=�F�u��y2�u.3�9~uV�/y  Y�;Fu9~u@���F@�t8t@����[_^]È�F�F�����F��%�   ��jh��<b  3�3�9u��;�u��D  �    VVVVV�����������+�u�lr  Y�u��u�u�����YY�E��E������	   �E��&b  ��u�r  YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�v  YP�  ��;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�Gv  P�/�  Y��Y��3�^]�jh8��a  3��}�}�j�V  Y�}�3��u�;5`+��   �@��98t^� �@�tVPV�q  YY3�B�U��@���H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u�@�4�V�q  YY��E������   �}�E�t�E��`  �j�{T  Y�jh`��@`  3�9uu	V����Y�'�u�p  Y�u��u����Y�E��E������	   �E��I`  ��u��p  Y�j�����Y�jh����_  3ۉ]�3��u;���;�u �B  �    SSSSS�}���������   �E��t	;�t��@u�;�t��@u�}�G�=���v뷋}����uV��o  Y�]�V����V�F  YY�f�����N�Et���Fj_�-�E;�u W�,  Y;�u�@�M����N  �	��   �N�~�F��^�E������	   �E��B_  ��u��o  YË�U���SVW3�9}t$9}t�u;�u�A  WWWWW�    ������3�_^[�ËM;�tڃ��3��u9Ew͋}�}�F  �M��}��t�F�E���E�   ����   �N��  t/�F��t(��   ��;�r��W�u��6�  )~>��+�}��O;]�rO��tV�S���Y��u}�}� ��t	3ҋ��u�+�W�u�V�s  YP�"|  �����ta��;�w��M�+�;�rP�}��)�E�� VP�s  YY���t)�E��FK�E����E�   ���A����E������N ��+�3��u������N �E���jh���]  3�9ut)9ut$3�9u��;�u �,@  �    VVVVV������3��]  ��u�m  Y�u��u�u�u�u�=������E��E������   �E����u��m  YË�U��W3�9}u��?  WWWWW�    ����������AV�u;�u�?  WWWWW�    �����������u��  Y�ȉ#ʃ���V;�t3�^_]Ë�U��V�u�F��u�P?  �    ����g���}�FuV�c�  E�e YV�����FY��y����F��t�t�   u�F   �u�uV�<q  YP�@�  3Ƀ������I��^]�jh���
\  3�3�9u��;�u�>  �    VVVVV����������>�};�t
��t��u��u�)l  Y�u�W�u�u�������E��E������	   �E���[  ��u�il  YË�U��V3�9uu�D>  VVVVV�    �0����������E;�t�V�p�0�u耂  ��^]Ë�U��SV�uW3����;�u��=  WWWWW�    ���������B�F�t7V�:���V����z  V�p  P��  ����}�����F;�t
P�&���Y�~�~��_^[]�jh����Z  �M��3��u3�;���;�u�u=  �    WWWWW�a����������F@t�~�E���Z  �V��j  Y�}�V�*���Y�E��E������   �ՋuV�1k  YË�U���u�T���u�H��3���tP�=  Y���]�3�]Ë�U��� WV�:  3�Y;�u��<  WWWWW�    ����������49}t޹����E�I   �u�u��M�;�w�E��u�E��u�uP�U��_�Ë�U��V�u�EPj �uhp��z�����^]Ë�U��Q�e� S�]��u3��   W��ru�{���vn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9}�r��?�@��I��F�@��I��<�@��I��2�@��I��(�M�E����t:u@A�E�9]�r�3�_[��� �	+����U��j
j �u�h�  ��]��5d�5  Y��t��j�u�  jj �g  ���H  ��U��EVW��u|P�oK  Y��u3��  �P9  ��u�K  ����  �\���+�֝  �L�j  ��}��5  ����  ��| 耚  ��|j �Q�  Y��u�H�   ��l  ��3�;�u19=H~��H9=�u���  9}u{�l  �g5  ��J  �j��uY�"5  h  j��  ��YY;��6���V�5(��5��}4  Y�Ѕ�tWV�[5  YY�X��N���V�����Y�������uW��7  Y3�@_^]� jh ��\W  ����]3�@�E��u9H��   �e� ;�t��u.����tWVS�ЉE�}� ��   WVS�r����E����   WVS謆���E��u$��u WPS蘆��Wj S�B�������tWj S�Ѕ�t��u&WVS�"�����u!E�}� t����tWVS�ЉE��E������E���E��	PQ��  YYËe��E�����3��V  Ë�U��}u��  �u�M�U�����Y]� ��������������̃= ��  ���\$�D$%�  =�  u�<$f�$f��f���d$�ޡ  � �~D$f( �f(�f(�fs�4f~�fT0�f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$螞  ���D$��~D$f��f(�f��=�  |!=2  �fT��\�f�L$�D$����f� �fV �fT�f�\$�D$���������������̃=�+ t-U�������$�,$�Ã=�+ t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$��jh ��YT  �e� �u;5l+w"j�JI  Y�e� V�QQ  Y�E��E������	   �E��eT  �j�EH  YË�U��V�u�����   SW�=`��=� u�`�  j讏  h�   蚓  YY�|+��u��t���3�@P���uV�S���Y��u��uF�����Vj �5��׋؅�u.j^9�t�u�D�  Y��t�u�{����76  �0�06  �0_��[�V��  Y�6  �    3�^]�������������U��WV�u�M�}�����;�v;���  ��   r�=�+ tWV����;�^_u^_]��D  ��   u������r*��$��0��Ǻ   ��r����$�0�$�1��$��0�0D0h0#ъ��F�G�F���G������r���$��0�I #ъ��F���G������r���$��0�#ъ���������r���$��0�I �0�0�0�0�0�0�0�0�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��0��111,1�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��2�����$�@2�I �Ǻ   ��r��+��$��1�$��2��1�1�1�F#шG��������r�����$��2�I �F#шG�F���G������r�����$��2��F#шG�F�G�F���G�������V�������$��2�I D2L2T2\2d2l2t2�2�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��2���2�2�2�2�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U��QSVW�5�,  �5���}��,  ��YY;���   ��+ߍC��rwW�Q�  ���CY;�sH�   ;�s���;�rP�u���  YY��u�G;�r@P�u���  YY��t1��P�4��+  Y��u�+  ���V�+  Y��EY�3�_^[�Ë�Vjj �G  ��V�h+  ������ujX^Ã& 3�^�jh@���N  贎  �e� �u�����Y�E��E������	   �E�� O  �蓎  Ë�U���u���������YH]�������������̺���a�  ����ܜ  �Ƀ=@t����$�  �����z�����������������̃��$�m�  �   ��ÍT$��  R��<$�D$tQf�<$t�Ю  �   �u���=< �C�  �   ����@�  �  �u,��� u%�|$ u��襮  �"��� u�|$ u�%   �t����-��   �=< ��  �   �����  ZË�U����\�3ŉE�SV3�W��9\u8SS3�GWh@�h   S�p���t�=\��H���xu
�\   9]~"�M�EI8t@;�u�����E+�H;E}@�E�\����  ;���  ����  �]�9] u��@�E �5l�3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�/  ��;�t� ��  �P�r���Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5p�SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w��.  ��;�tj���  ���P����Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�p���t"SS9]uSS��u�u�u�VS�u �h��E�V�����Y�u�������E�Y�Y  �]�]�9]u��@�E9] u��@�E �u�`�  Y�E���u3��!  ;E ��   SS�MQ�uP�u �~�  ���E�;�tԋ5d�SS�uP�u�u�։E�;�u3��   ~=���w8��=   w��-  ��;�t����  ���P����Y;�t	� ��  �����3�;�t��u�SW�n������u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��ͬ  ���u������#u�W�����Y��u�u�u�u�u�u�d���9]�t	�u��\���Y�E�;�t9EtP�I���Y�ƍe�_^[�M�3������Ë�U����u�M������u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap�����(  �ȋAl;�t�0��Qpu�  ���   Ë�U����u�M������E����   ~�E�Pj�u��  ������   �M�H���}� t�M��ap��Ë�U��=d u�E���A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u� �  ������   �M�H���}� t�M��ap��Ë�U��=d u�E���A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u聬  ������   �M�H���}� t�M��ap��Ë�U��=d u�E���A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Ph�   �u���  ������   �M�H%�   �}� t�M��ap��Ë�U��=d u�E���A%�   ]�j �u�~���YY]Ë�U����u�M������E����   ~�E�Pj�u�|�  ������   �M�H���}� t�M��ap��Ë�U��=d u�E���A��]�j �u����YY]Ë�U���L�\�3ŉE�S3�V�uW�]ԉ]�]��]؉]܉u��]�9^�  �F9u P�F0h  P�E�SP�X�  ������  j�  j��  W�E��  jW�E��  jW�E��  jh  �E��  ��$�E�9]��|  9]��s  ;��k  9]��b  9]��Y  �Eԉ3��M܈@=   |�E�P�v�t����/  �}��%  �E���E�~-8]�t(�E�:�t�x�����M�� �G;�~�@@8X�uۋE�SS�v   Ph   �u܉E�jS�A�  �� ����  �M��E�S�v��   W���   QW@Ph   �vS������$����  �E�S�v�   WP�E�W@Ph   �vS�U�����$���`  �E�}����   3҃}�f��U؉Mč��   �_�Z��M����   �MȈ~S8]�tN�M�M�:�tB�I���;ʉM�'��H   ��M��E� �  f�AA�M̋M��	9M�~�M�AA�M�8Y�u�h�   ��   QP�]���j��   PW�N����E�j��   QP�<������   ��$;�tKP����u@���   -�   P�������   ��   +�P�������   +�P�u������   �j������E��    ���   �E����   �Eĉ��   �E����   �Eȉ��   �EЉ��   �u��#���Y���m�u������u������u������u������3ۃ�C�ˍ��   �;�tP������   ǆ�   H�ǆ�   Чǆ�   P�ǆ�      3��M�_^3�[�&������|"  �ȋAl;�t�0��Qpu�r  �@��V"  �ȋAl;�t�0��Qpu�L  ��Ë�U��VW3��u�������Y��u'9`vV�����  ;`v��������uʋ�_^]Ë�U��VW3�j �u�u蕩  ������u'9`vV�����  ;`v��������uË�_^]Ë�U��VW3��u�u�i�  ��YY��u,9Et'9`vV�����  ;`v��������u���_^]Ë�U��VW3��u�u�u�3�  ������u,9Et'9`vV�����  ;`v��������u���_^]��̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U���(  �\�3ŉE����Vtj
��|  Y��  ��tj��  Y�����   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P�f�������������(�����0���j ǅ����  @��������,����<���(���P�8�j��  ̋�U��M����U#U��#�ʉ��]�Pd�5    �D$+d$SVW�(��\�3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(��\�3�P�e��u��E������E�d�    ËM�d�    Y__^[��]QË�U��SV�u���   3�W;�to= th���   ;�t^9uZ���   ;�t9uP�������   �0�  YY���   ;�t9uP�������   � �  YY���   �j������   �_���YY���   ;�tD9u@���   -�   P�>������   ��   +�P�+������   +�P�������   ���������   �=@t9��   uP�m�  �7�����YY�~P�E   ��8�t�;�t9uP�����Y9_�t�G;�t9uP����Y���Mu�V����Y_^[]Ë�U��SV�5�W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�8�t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5�W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�8�t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�V���t��t;�tWj6Y���  P����Y_^Å�t7��t3V�0;�t(W�8����Y��tV�����> Yu��@�tV�3���Y��^�3��jh`��<  ��  ��0��Fpt"�~l t��  �pl��uj ��{  Y����<  �j�1  Y�e� �Fl�=��i����E��E������   ��j�0  Y�u�á��H���H�����   �����   �����   �0���   ������   �4�3�Ë�U��SW�}3�;�~,V�u���6�u�u�
�  ����tSSSSS�c�����Ou�^_[]Ë�U��SVW�}h�   3�SW�����u�����u3���   <.u4�F8t-jP���   jP�m�  ����tSSSSS����������   ��hX�V�]���  ;��   �} �<0�u��@��   ��.��   PVj@�u�;�}u��@sw��_trP�EVj@��@��}u`��s[��t��,uRP�EVj��P�ֳ  ����t3�PPPPP�f�������,�'����������E�whX�V�X�  ��YY�X������_^[]Ë�U��SV�uV�u�u�������3ۅ�tSSSSS�������F@8tPh\�j�u�u�Q��������   8^[tPh�j�u�u�/�����]Ë�U���S3�ChU  �]������Y�E���U  W�x� ��]��^�CH�0�E�hd��5��jhQ  W������E���E��E���h`�hQ  W��  ����t3�PPPPP�;������sX�E��0�  YY��t�e� �E��E��E����0�CH�0�E�E�hd��0jhQ  W�Z������}�̪|��}� uI�FP����tP�Ӆ�u	�vP�n���Y�FT��tP�Ӆ�u	�vT�W���Y�E�fT �fL �FP�~H���N�u��9����FP�=�3�Y;�tP�ׅ�u	�vP����Y�FT;�tP�ׅ�u	�vT����Y�Fh�^T�^L�^P�^H_[�Ë�U���   �\�3ŉE��ESV�uW�}��d����E��\�����`����  �   �H(��T����H,�X �   ��X�����h�������  ��d��� ��  �} ��  �>CuW�~ uQh���u��d����l�����3���tVVVVV������;�t3�f�f�Gf�G��`���;�t�0��d����G  V�������   Y��P���;�s,V��h����  YY����   V��X����  YY����   ��L��� ��l���VP����YY����   ��l���PSP�ɶ  ������   �C��T������l���PW��h����������> t
��P���;�r��L������@PVW��X�����  ����t3�VVVVV�������3�9�\���tjS��\���������9�`���tj��T�����`�����������h����u��d�����������tVVVVV�0�������h����3��M�_^3�[�B����Ë�U����  �\�3ŉE�SW���  �u����h���P��P���Ph�   ��x���PS���  ��������u3��  �E���0�sH��x���P��
  YY���x  ��x���P������P��t��������YY��p�����t��CH�M��\����D���k���l���� ��X����1jP��d�����<���P�_����F��x���Q��t�����L�����p��������QP���������t3�PPPPP���������p�����l������CH��P����j��P���P��d�����������}��   ��h�����t��� �F�G$�O ��d����ǋV;t6���t������d�����D����P�H��D�������t�����d���|��"��t�����t�ǋ��P�W���d����H��t���uhj�v��x����vPjhتjj ��  �� ��t93���  f!�Ex���@��r�h�   �5����x���P裵  �����@�G��g �F��G���   �}u	��h����F�Ek�V����Y��t1��\�����p����CH�;�����X���Y��l������L����F������\���8�t-�E�����<0�7����u�7������sT������cL YY�M��p��������    �1�CH�M�_3�[�@����Ë�U���   �\�3ŉE��ESV3ۋ�W��h���;�t;�tP�����Y��  ���D0H��  ǅp���   ��t���;���  �9L�0  �yC�&  �y_�  ��hh�W���  ��YY����   +ǉ�p�����   �;;��   ǅl���   ������p���PW�6��������u�6�����Y9�p���t��l�������̪~�Ch`�S�+�  ��3�YY;�u	�;;��   ��l���QWS��x���h�   P�B�  ����tVVVVV���������l�����h�����x���Ƅ=x��� ����Y��t��t�����? t
G�? � ���3�9�t�����   ��h����u3��vSSSh�   ��x���PQ�"�����;�tZ�~H��t3�7��x���P�  YY��tS��x����%���Y��u!�p������t���C����~�3�9�p���u9�t���t�D����M�_^3�[�%�����jh���R1  3ۉ]��}v�  �    SSSSS�������3��,  �E  ���u��N����Np�]�jh�   �8���YY���}�;���   j��%  Y�E�   �Nl�������]��   �u�M���P���Y�E�;���   9]th8��u�  YY��t
�d   j�%  Y�E�   �^l���y���W����Y�Fpu2�0�u)�;���W���j����Ph�������������e� �   �-�}܋u�3�j�V$  YËu�j�J$  Y��W�K���W�m���YY�E������   �E��<0  Ëu�fp��jh����/  3��u�3��];���;�u�  �    VVVVV�{�����3��{3��};���;�t�3�f97��;�t��h�  �E;�u�M  �    �ɉu�f93u �8  �    j��E�Ph\��i�  ���P�uWS�m�  ���E��E������	   �E��x/  ��u� @  YË�U���SV�u3ۉ]�;�t9]u3��{  v3�f�W�};�u�  SSSSS�    �������<  �u�M��v����E�;���   9XuH9]v�M��9f�f�8tAFF�M�;Mr�8]�t�E�`p��E���   8]�t�E�`p�����   �uVj�W�=l�j	�p��;���   �H���zt�  � *   3�f��   �E�u�E�;�t'��M�:�t�M���QP�w�  YY��tF8t!F9]�u��u+u�u�E�V�uj�p��;�uT�  �M� *   3�f��-9Xu	W�����Y�1SSj�Wj	�p�l�;�u�u  � *   8]�t�E�`p�����H8]�t�M�ap�_^[�Ë�U���SV�u3ۉ]�;�u9]t*�9]w�%  j^SSSSS�0����������   3�f�W�};�t��u�M��Զ���E;Ev�E=���v	��  j�P�M�QP�uV����������u;�t3�f��  � 8]�tk�M�ap��b@;�tH;Ev<�}�t,3�f��  j"^SSSSS�0�v�����8]�t�E�`p����&�E�E�P   3�f�LF�;�t�8]�t�E�`p��E�_^[�Ë�U��j �u�u�u�u�u�������]�������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[�jh���v+  j�v   Y�e� �u�N��t/�l�h�E��t9u,�H�JP����Y�v�y���Y�f �E������
   �e+  Ë���j�A  Y��̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�"���3��ȋ��~�~�~����~��������F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �\�3ŉE�SW������P�v�t��   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R�_�����C�C��u�j �v�������vPW������Pjj ��  3�S�v������WPW������PW�vS�C�����DS�v������WPW������Ph   �vS������$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[�)�����jh���V(  �s  ���0��Gpt�l t�wh��uj �g  Y���n(  �j�(  Y�e� �wh�u�;58�t6��tV����u���tV�4���Y�8��Gh�58��u�V���E������   뎋u�j��  YË�U���S3�S�M��Q����p���u�p   �|�8]�tE�M��ap��<���u�p   �x��ۃ��u�E��@�p   ��8]�t�E��`p���[�Ë�U��� �\�3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�@���   �E��0=�   r����  �p  ����  �d  ��P������R  �E�PW�t����3  h  �CVP����3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�8����M��k�0�u���P��u��*�F��t(�>����E���<�D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C��D�Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95p�X�������M�_^3�[�$�����jh��Q%  �M���j  ���}�������_h�u�u����E;C�W  h   �
���Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh����u�Fh=�tP����Y�^hS�=����Fp��   �0���   j�  Y�e� �C���C���C��3��E��}f�LCf�Et@��3��E�=  }�L��0�@��3��E�=   }��  ��8�@���58�����u�8�=�tP�W���Y�8�S���E������   �0j�"  Y��%���u ���tS�!���Y�  �    ��e� �E��	$  Ã= uj��V���Y�   3�Ë�U��V�5,��5���օ�t!�(����tP�5,����Ѕ�t���  �'�|�V�����uV�b  Y��thl�P�����t�u�ЉE�E^]�j ����YË�U��V�5,��5���օ�t!�(����tP�5,����Ѕ�t���  �'�|�V�����uV�b  Y��th��P�����t�u�ЉE�E^]����� ��V�5,��������u�5��e���Y��V�5,������^á(����tP�5��;���Y�Ѓ(���,����tP����,���  jh8��2"  �|�V�����uV�Ua  Y�E�u�F\0�3�G�~��t$hl�P����Ӊ��  h���u��Ӊ��  �~pƆ�   CƆK  C�Fh�j��  Y�e� �vh���E������>   j�  Y�}��E�Fl��u���Fl�vl�+���Y�E������   �!  �3�G�uj�  Y�j�  YË�VW�H��5(��������Ћ���uNh  j�^�����YY��t:V�5(��5������Y�Ѕ�tj V�����YY�X��N���	V�0���Y3�W���_��^Ë�V��������uj�2`  Y��^�jh`��   �u����   �F$��tP����Y�F,��tP�ն��Y�F4��tP�Ƕ��Y�F<��tP蹶��Y�F@��tP諶��Y�FD��tP蝶��Y�FH��tP菶��Y�F\=0�tP�~���Yj�:  Y�e� �~h��tW����u���tW�Q���Y�E������W   j�  Y�E�   �~l��t#W����Y;=�t��@�t�? uW�)���Y�E������   V�����Y��  � �uj��  YËuj��  YË�U��=(��tK�} u'V�5,��5���օ�t�5(��5,����ЉE^j �5(��5�����Y���u�x����,����t	j P���]Ë�VW�|�V�����uV�F^  Y�����^  �5��hȫW��h��W����h��W����h��W���փ=� �5����t�=� t�=� t��u$����������`�5�������,������   �5�P�օ���   �S`  �5������5��������5��������5����u��������  ��teh�a�5������Y�У(����tHh  j������YY��t4V�5(��5�����Y�Ѕ�tj V�y���YY�X��N��3�@��$���3�_^Ë�U��3�9Ev�M�9 t@A;Er�]Ë�U��E3�;�0�tA��-r�H��wjX]Ë�4�]�D���jY;��#���]��������u���Ã���������u���Ã�Ë�U��V������MQ�����Y�������0^]���Q�L$+ȃ����Y銺  Q�L$+ȃ����Y�t�  ��U���(  ���������5��=�f��f��f��f��f�%�f�-�����E ���E���E���������  ������	 ���   �\��������`��������@��j��  Yj �<�hԫ�8��= uj�  Yh	 ��4�P�0���U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh����  �e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E���  Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[��������+3�Ë�U���V�u�M�謣���u�P��  ��e�F�P������Yu��P���  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M��9����E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�:�  �M��E��M��H��EP�ɸ  �E�M����Ë�U��j �u�u�u������]Ë�V����tV����@PV�V�r�����^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M��������3�;�u+�	���j_VVVVV�8��������}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�����j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]hܫSV�ޣ����3ۅ�tSSSSS�������N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F�t�90uj�APQ�������}� t�E��`p�3�_^[�Ë�U���,�\�3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�ܸ  3ۃ�;�u�~���SSSSS�0�n��������o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q���  ��;�t���u�E�SP�u��V�u��������M�_^3�[�����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   芟��9}}�}�u;�u+����j^WWWWW�0聫�����}� t�E�`p����  9}vЋE��� 9Ew	�V���j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�߲  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� 觷  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �S�  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�[�����u�E�8 u���} �4����$�p���WF�߶  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP躵  0�F�U�����;�u��|��drj jdRP蔵  0��U�F����;�u��|��
rj j
RP�n�  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N������u-�3���j^�03�PPPPP�������}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V蕞�����}� t�E��`p�3�_^[�Ë�U���,�\�3ŉE��ESVW�}j^V�M�Q�M�Q�p�0肳  3ۃ�;�u�$���SSSSS�0���������Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P谱  ��;�t���u�E�SV�u���`������M�_^3�[誝���Ë�U���0�\�3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�ǲ  3ۃ�;�u�i���SSSSS�8�Y��������   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW���  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[谜���Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3������6������Y���(r�_^Ë�Vh   h   3�V���  ����tVVVVV萣����^Ë�U������]����]��E��u��M��m��]����]�����z3�@��3���h������th��P�����tj �������U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]Ã%�+ Ë�U��3�9Ej ��h   P�������u]�3�@�|+]Ã=|+uWS3�9d+W�=L�~3V�5h+��h �  j �v�����6j �5��׃�C;d+|�^�5h+j �5���_[�5�����%� Ë�VW3����<���u�����8h�  �0���{�  YY��tF��$|�3�@_^Ã$��� 3����S�$�V���W�>��t�~tW��W�H����& Y����� |ܾ��_���t	�~uP�Ӄ���� |�^[Ë�U��E�4����,�]�jh���  3�G�}�3�9�u�I  j�[G  h�   �GK  YY�u�4���9t���nj�\���Y��;�u�(����    3��Qj
�Y   Y�]�9u,h�  W�r�  YY��uW�v���Y������    �]���>�W�[���Y�E������	   �E��H  �j
�(���YË�U��EV�4����> uP�"���Y��uj�;J  Y�6�(�^]Ë�U��d+�h+k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �8����   �x+�5��h @  ��H� �  SQ�֋x+�8�   ���	P�8�@�x+����    �8�@�HC�8�H�yC u	�`��8�x�ueSj �p�֡8�pj �5��L��d+�8k��h++ȍL�Q�HQP蕕���E���d+;8v�m�h+�p+�E�8�=x+[_^�át+V�5d+W3�;�u4��k�P�5h+W�5����;�u3��x�t+�5d+�h+k�5h+h�A  j�5��`��F;�t�jh    h   W����F;�u�vW�5��L�뛃N��>�~�d+�F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�����u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U����d+�Mk�h+������M���SI�� VW}�����M���������3���U��p+����S�;#U�#��u
���];�r�;�u�h+��S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1�h+�	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t�p+�C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;8u�M�;x+u�%8 �M���B_^[����h �d�5    �D$�l$�l$+�SVW�\�1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s35\�W��E� �E�   �{���t�N�38�,����N�F�38�����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t����  �E���|@G�E��؃��u΀}� t$����t�N�38詋���N�V�3:虋���E�_^[��]��E�    �ɋM�9csm�u)�= � t h ��ӣ  ����t�UjR� ����M賛  �E9Xth\�W�Ӌ�趛  �E�M��H����t�N�38�����N�V�3:�����E��H���I�  �����9S�R���h\�W���a�  ������U��V�EP��蘏���(���^]� �(��0�����U��V���(������EtV�u��Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR����YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =MOC�t=csm�u+�h������    ��  �W������    ~�I����   �3�]�jh�������}�]��   �s��s�u������   � �e� ;ute���~;w|��  �����Oȋ1�u��E�   �y t�sh  S�O�t��  �e� ��u��-���YËe�e� �}�]�u��u���E������   ;ut�V  �s����Ë]�u��s������    ~�e����   �Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�'���3�A��  ���3��jh��������M��t*�9csm�u"�A��t�@��t�e� P�q�Ò���E�����������3�8E��Ëe��G
  ̋�U��M�V�uƃy |�Q�I�42���^]Ë�U�����u
�X
  �
  �e� �? �E� ~SSV�E�@�@��p��~3�E����E�M�q�P�GE�P�_�������u
K�������E��E��E�;|�^[�E���j�ό�����������    t��	  �e� �	  �M���q	  ������Mj j ���   謐���j,hh������ً}�u�]�e� �G��E��v�E�P�9���YY�E��������   �E��������   �E��������   �x����M���   �e� 3�@�E�E��u�uS�uW臔�����E�e� �o�E������Ëe��5�����   �u�}�~�   �O��O�^�e� �E�;Fsk�ËP;�~@;H;�F�L�QVj W�������e� �e� �u�E������E    �   �E��������E�맋}�u�E܉G��u�腓��Y�����Mԉ��   �����MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v����Y��t�uV�%���YY�jh������3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w觞  YY����   SV薞  YY����   �G��M��QP�����YY���   �}�E�p�tH�_�  YY����   SV�N�  YY����   �w�E�pV�(��������   ���t|��W�9Wu8��  YY��taSV��  YY��tT�w��W�E�p�_���YYPV�ׅ�����9�ڝ  YY��t)SV�͝  YY��t�w违  Y��t�j X��@�E���  �E������E��3�@Ëe��F  3�������jh�������E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS�>�����FP�w����YYP�vS�$����E������Z����3�@Ëe��  ̋�U��} t�uSV�u�V������}  �uuV��u �����7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP�l���]Ë�U��QQV�u�>  ���   W�������    t?�������   �0���9t+�>MOC�t#�u$�u �u�u�u�uV����������   �}� u�  �u�E�P�E�PV�u W�N������E���;E�s[S;7|G;wB�G�O����H��t�y u*�X��@u"�u$�u�u j �u�u�u�u�����u���E��E���;E�r�[_^�Ë�U���,�MS�]�C=�   VW�E� �I��I����M�|;�|�]  �u�csm�9>��  �~� ��  �F;�t=!�t="���   �~ ��   �G������    ��  �5������   �u�'������   jV�E��  YY��u��  9>u&�~u �F;�t=!�t="�u�~ u�  ��������    t|��������   ������u3����   ����Y��uO3�9~�G�Lh� ��}����uF��;7|��	  j�u�d���YYh0��M��7���h���E�P�4����u�csm�9>��  �~�~  �F;�t=!�t="��e  �}� ��   �E�P�E�P�u��u W�&��������E�;E���   �E�9��   ;G|�G�E�G�E��~l�F�@�X� �E��~#�v�P�u�E����������u�M��9E���M�E��}� ��(�u$�]��u �E��u��u�u�uV�u�K����u���E����]����}�} t
jV�:���YY�}� ��   �%���=!���   �����   V����Y����   ���������������   � ����}$ �M���   Vu�u��u$�ˉ���uj�V�u�u�������v�����]�{ v&�} �)����u$�u �u�S�u�u�uV������� �������    t�T  _^[�Ë�U��V�u���6����(���^]� ��U��SVW�V�����   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������� 3�@_^[]�jh��O����l����@x��t�e� ���3�@Ëe��E������ӯ���h�����?����@|��t������jh(������5<�����Y��t�e� ���3�@Ëe��E������}����he��(���Y�<�������U���SQ�E���E��EU�u�M�m�詗  VW��_^��]�MU���   u�   Q臗  ]Y[�� � á`+Vj^��u�   �;�}�ƣ`+jP�y���YY�@��ujV�5`+�`���YY�@��ujX^�3ҹ ��@��� �����|�j�^3ҹ0W������@����������t;�t��u�1�� B���|�_3�^�迏���=� t��  �5@����YË�U��V�u� ;�r"���w��+�����Q�z����N �  Y�
�� V�(�^]Ë�U��E��}��P�M����E�H �  Y]ËE�� P�(�]Ë�U��E� ;�r=�w�`���+�����P�*���Y]Ã� P�,�]Ë�U��M���E}�`�����Q�����Y]Ã� P�,�]Ë�U��V�uW3�;�u�o���WWWWW�    �[�������   �F����   �@��   �t�� �F��   ���F�  u	V�  Y��F��v�vV�W  YP�ڛ  ���F;���   �����   �F�uOV�-  Y���t.V�!  Y���t"V�  ��V�<�@�  ��Y��Y����@$�<�u�N    �~   u�F�t�   u�F   ��N�A���������	F�~���_^]�jThH�����3��}��E�P�Đ�E�����j@j ^V虪��YY;��  �@�5 ��   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@�@��   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M���@��  ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9= |���= �e� ��~m�E����tV���tQ��tK�uQ�����t<�u���������4�@�E� ���Fh�  �FP�O�  YY����   �F�E�C�E�9}�|�3ۋ���5@����t���t�N��r�F���uj�X�
��H������P��������tC��t?W�����t4�>%�   ��u�N@�	��u�Nh�  �FP蹏  YY��t7�F�
�N@�����C���g����5 ���3��3�@Ëe��E������������Ë�VW�@�>��t1��   �� t
�GP�$����@   ;�r��6�G����& Y����@|�_^Ë�U��EV3�;�u����VVVVV�    菀���������@^]Ë�U��QV�uV�����E�FY��u�e���� 	   �N ����/  �@t�J���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,������� ;�t�������@;�u�u�Z�  Y��uV��   Y�F  W��   �F�>�H��N+�I;��N~WP�u�  ���E��M�� �F����y�M���t���t�����������@����@ tjSSQ軘  #����t%�F�M��3�GW�EP�u�  ���E�9}�t	�N �����E%�   _[^�Ë�U���@h   �4���Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U���  贆  �\�3ŉE��EV3���4�����8�����0���9uu3���  ;�u'�����0����VVVVV�    �w~��������  SW�}�����4�@�����ǊX$�����(�����'�����t��u0�M����u&�<���3��0� ���VVVVV�    �~�����C  �@ tjj j �u�Ė  ���u�W�  Y����  ��D���  �+����@l3�9H�������P��4�� ����А���`  3�9� ���t���P  �̐��4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P��  Y��t:��4���+�M3�@;���  j��@���SP蠙  �������  C��D����jS��@���P�|�  �������  3�PPj�M�Qj��@���QP�����C��D����h������\  j ��<���PV�E�P��(���� �4�Ȑ���)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4�Ȑ����  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@���艖  Yf;�@����h  ��8����� ��� t)jXP��@����\�  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4�Ȑ���B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4�Ȑ���b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �h���;���   j ��,���P��+�P��5����P��(���� �4�Ȑ��t�,���;����H���@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0�Ȑ��t��,�����@��� ��8�����H���@�����8��� ul��@��� t-j^9�@���u����� 	   �����0�?��@�������Y�1��(�����D@t��4����8u3��$������    ������  ������8���+�0���_[�M�3�^�n����jhh�������E���u�����  ����� 	   ����   3�;�|; r!�v����8�\���� 	   WWWWW�Hw�����ɋ�����@��������L1��t�P�g�  Y�}���D0t�u�u�u�.������E�������� 	   �����8�M���E������	   �E��T�����u豕  Y�jh��������E���u����� 	   ����   3�;�|; r����� 	   SSSSS�{v�����Ћ����<�@��������L��t�P蚔  Y�]���Dt1�u��  YP�Ԑ��u�H��E���]�9]�t�.����M������ 	   �M���E������	   �E��s�����u�Д  YË�U��V�u�F��t�t�v�Jv���f����3�Y��F�F^]Ë�U��   �}  �\�3ŉE�SV�uWV�������3�9FY������}�FjPPS�ʎ  ������������������|��s
������  ������@��������� ��ÊH$����F  ������u�F�������+�ʋǋ��  ��V��+��V���������Z  �������  3�9P0�  �����9Vu�������������<  R�p,�p(���������  ��������� Ã���;p(�0���;x,�'���j ������Qh   ������Q�0�ؐ������j ������������������蘍  ����������������������������;��������������t7������K;�s+���u�J�;�s�H�9
u�������P�@��uЍ�����+�3����L  �@�t�V��:
u������B;�r������������u�������  ��x������    �$����F��   �V��u!�������   +N��@�����   jj j ������蕌  ��;�����u$;�����u�F�8��8
uG@;�r��F    �Yj �������������������M�  �����������������   ;�w�N��t
����   t�~������� �DtG������u��)����������� ������uѭ����������3������������M�_^3�[�mi����jh�������u�����Y�e� �u����Y�E��U��E������   �E��U�������u�4���YË�U��V�uV��  Y���u����� 	   ����MW�uj �uP�ܐ�����u�H��3���tP�����Y����������@�����D0� ���_^]�jh��������E���u覾���  苾��� 	   ����   3�;�|; r!�}����8�c���� 	   WWWWW�Oq�����ɋ�����@��������L1��t�P�n�  Y�}���D0t�u�u�u��������E��� ���� 	   �����8�M���E������	   �E��[�����u踏  YË�U���SW�}3�;�u 踽��SSSSS�    �p��������f  W�����9_Y�E�}�_jSP�������;ÉE�|ӋW��  u+G�.  ��OV��+�u���tA�U��u�����@�����D2�t��;�s���:
u�E�3�B;�r�9]�u�E���   ��x��	����    �   �G��   �W;�u�]��   �]��u�+��������@�E����D0�tyjj �u�������;E�u �G�M��	�8
u�E@;�r��G    �@j �u��u����������}����:�   9Ew�O��t��   t�G�E��D0t�E�E)E��E�M��^_[�Ë�U��V�u�FW��ty�}��t
��t��uh���F��uV�I���EYU3�V�Vw���FY��y����F��t�t�   u�F   W�u�uV����YP��  #����t3��褻���    ���_^]�jh��������u�!���Y�e� �u�u�u�u�:������E��E������	   �E��������u�[���YË�U��V�uWV��  Y���tP�@��u	���   u��u�@Dtj�܋  j���Ӌ  YY;�tV�ǋ  YP� ���u
�H����3�V�#�  ������@����Y�D0 ��tW�޺��Y����3�_^]�jh�������E���u覺���  苺��� 	   ����   3�;�|; r!�}����8�c���� 	   WWWWW�Om�����ɋ�����@��������L1��t�P�n�  Y�}���D0t�u�����Y�E������� 	   �M���E������	   �E��j�����u�ǋ  YË�U��9EuF�jP;Mu+�1���YY���u3�]ËE�    �6�u�7螃�����Q蟔������tՉ�&3�@]Ë�U���EP耎�����EYu��߃�]��Jx	�
�A�
�R�����YË�U��}�t]�Cs��]Ë�U��S�U�������؃��t��P�+���Y��u��[]Ë�U����  �\�3ŉE��M�EV3�W�}�������|�����d�����T���ǅ$���^  ��0����������x���;�u 趸��VVVVV�    �k��������5  ;�t��@@SuzP�����Y�����t���t�ȃ��������@����A$u&���t���t�ȃ������@����@$�t �1���VVVVV�    �k��������  �u�������^���ƅc��� ��t�����<������k  ��d�����P����Y��t0��t���VV��t�������YP�k���YYG�P轍��Y��u��  �<%�1  8G�  3���@���ƅ/��� ��X�����L�����l���ƅa��� ƅ`��� ƅj��� ƅS��� ƅb��� ƅs��� ƅk�����(���G���P�6���Y��t��l�����L���k�
�DЉ�l�����   ��N��   ��   ��*tp��F��   ��It��Lut��k����   �O��6u�G�84u��(�������4�����8����m��3u�G�82u���\��dtW��itR��otM��xtH��Xu�A��j����9��ht(��lt��wt��S����"�G�8lt���k�����s������k�����s�����S��� �������j��� ��H���u������0�������������3�2ۉ�D���8�s���u�<Stƅs����<Cuƅs������ ��\�����ntJ��ct��{t��d�����t����}���Y���d�����t����@�����x��������  ��D�����H�����L�����t��l��� ��  ��\�����o�r  �  ��c�
  jdZ;���  �z  ��g~E��it!��n�g  ��j��� ��t����f
  �
  ��\�����x���-�4  ƅ`����1  3ۃ�x���-u��T���� -C�	��x���+u��l�����d�����t����^�����x�����L��� u��l������x����k��l�����l�����tf��x�����T�����X������0���P��|���PCS��T�����$�������������
  ��d�����t����������x�����P�=���Y��u���������   � � ��a���:�x�����   ��l�����l�������   ��d�����t���������T�����x�����a������0���P��|���PCS��T�����$��������������	  ��x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$����{���������	  ��d�����t����������x�����P�6���Y��u���X��� �_  ��x���et��x���E�I  ��l�����l������5  ��T����e��0���P��|���PCS��T�����$��������������  ��d�����t����D�����x�����-u,��T����-��0���P��|���PCS����������  �	��x���+u/��l�����l�����u!�l������d�����t����������x�����x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$������������  ��d�����t����j�����x�����P�ʆ��Y��u���d�����t�����x����U�����X��� YY��  ��j��� ��  ��T�����<��������QP��D���� ��k���HP�5���j���Y�Ѓ��  ��u��l���ǅL���   ��s��� ~ƅb�����d�����t���W��x�����@�������YY��L��� t��l�����l������3  ��t������x�����x�������  ��\���ctN��\���su��	|	����  �� u2��\���{��  ��a���3ҋȃ�B������L�3˅���  ��j��� ��  ��b��� �~  �� �����P�#k  Y��t��t������������!��������P�����ǅ���?   ���   �� ���P�����P�~  f�������f�FF�  ��p��  �������HH�{  ���������t3�;�x�����  ��c�����j��� �  �����������  ��s��� ~ƅb���G�?^��u
�wƅa����j �E�j P�Y�����>]u	�]F�E� �f��/����^F<-uB��t>���]t7F:�s�����:�w"*������Ћσ��ǳ�����D�GJu�2���ȊЋ��������D��<]u����  ��H�����D���������x���+u'��l���u��t����d�����t����C�����x���j0^9�x����x  ��d�����t���������x���<xtX<XtT��\���xǅX���   t"��L��� t
��l���u��ǅ\���o   �$  ��d�����t���P�����YY��x����  ��d�����t���������L��� ��x���t��l�����l���}��ǅ\���x   ��   �F��D����������@���������t���WP�j���YY9�@�����  ��j��� �  ��<�����\���c��  ��b��� t��D���3�f���  ��D����  ��  ƅk�����x���-u	ƅ`����	��x���+u'��l���u��t����d�����t���������x�����(��� �J  ���  ��\���xte��\���pt\��x���P����Y����   ��\���ou"��x���8��   ��4�����8��������Rj j
��8�����4����,[�������7��x���P����Y��tr��4�����8�����x������������Y��x�����x�����X�����Й����L��� ��4�����8���t��l���t5��d�����t���������x���������d�����t�����x�������YY��`��� ��@�����   ��4�����8����؃� �ى�4�����8�����   ��@�������   ��\���xt;��\���pt2��x���P血��Y����   ��\���ou��x���8}n���,k�
�'��x���P����Y��tR��x����������Y��x�����X�����L��� ��x����|�t��l���t5��d�����t���������x����X�����d�����t�����x�������YY��`��� t�߃�\���Fu��X��� ��X��� �  ��j��� u8��<�����D�����(��� t��4������8����F���k��� t�>�f�>��H�����c���G��H����`<%u
�G�8%u����t�������������G��x�����H���;�ul��P�e  Y��t!��t�����������G��H���;�uG��t�����x����u�?%uD��H����xnu8������	����*��d�����x�������YY�VS��VP����VS�y�������0���u��T����2]��Y��x����u*��<�����u8�c���u�������� t%������ap������� t
������`p���<���[�M�_3�^�ZS���Ë�U���VW�u�M��%P���E�u3�;�t�0;�u,�,���WWWWW�    �\�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�4*  �M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&苧���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9duh ��P������]Ë�U��QQS�]VW3�3��}�;��t	G�}���r���w  j�q|  Y���4  j�`|  Y��u�=X�  ���   �A  h��  S�HW�P������tVVVVV�FX����h  �aVj �e �����u&hбh�  V��O������t3�PPPPP�X����V老��@Y��<v8V�s�����;�j�\ẖ+�QP�/<  ����t3�VVVVV�W�����3�hȱSW�B;  ����tVVVVV�W�����E��4��SW�;  ����tVVVVV�vW����h  h��W��y  ���2j������;�t$���tj �E�P�4���6辀��YP�6S�Ȑ_^[��j��z  Y��tj��z  Y��u�=Xuh�   �)���h�   ����YYË�U���   �\�3ŉE��ESV�u3ۃ}W��t�����l�����   Sh�   ��|�����Q�u��x����uP�*|  ����;�uj�H���z��   SSS�u�u��t�����{  ����p���;�t_3�FVP��~����YY;�tMS��p�����x���W�u�u��t�����{  ����;�tjV�~��YY��l����;�u!9�x���tW�W��Y����M�_^3�[�N���ÍN�QWVP�>:  ����tSSSSS��U����9�x���tW�iW��Y3��9]u�Sj�\W�u�uP��y  ����t�����P�x��Y��tɊ�
���,0GG��d�|�뱋�U��E�d]Ë�U��W��  W���u������  ��`�  w��t�_]Ë�U��������u�L����5��P���h�   �Ѓ�]Ë�U��h������th�P�����t�u��]Ë�U���u�����Y�u���j�+���Y�j�H���YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=�� th����d  Y��t
�u���Y�n���h��hx�����YY��uBh����p���\��$t��c����= Yth�d  Y��tj jj �3�]�jh(��G���j�G���Y�e� 3�C9���   ���E���} ��   �5�ߛ��Y���}؅�tx�5�ʛ��Y���u܉}�u����u�;�rW覛��9t�;�rJ�6蠛����萛������5芛�����5�}�����9}�u9E�t�}�}؉E����u܋}��h������_���Yh������O���Y�E������   �} u(��j�u���Y�u�����3�C�} tj�\���Y��m���Ë�U��j j�u�������]�jj j ������Ë�V�ǚ����V�
  V�b  V�pR��V�
���V�Cx  V�e(  V�(K��V�����h��������$��^Ã= u����V�5LW3���u����   <=tGV�{��Y�t���u�jGW�z����YY�=x��tˋ5LS�BV�t{����C�>=Yt1jS�uz��YY���tNVSP�I������t3�PPPPP�Q�������> u��5L�KS���%L �' �   3�Y[_^��5x�%S���%x ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�Gw  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�bv  Y��t��M�E�F��M��E���?v  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9u�_���h  ��VS�������+�5�;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�w����Y;�t)�U��E�P�WV�}�������E���H�l�5p3�����_^[�Ë�U�졨��SV�5��W3�3�;�u.�֋�;�t��   �#�H���xu
jX���������   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5h�SSS+�S��@PWSS�E��։E�;�t/P��v��Y�E�;�t!SS�u�P�u�WSS�օ�u�u�� P��Y�]��]�W�����\��t;�u�����;��r���8t
@8u�@8u�+�@P�E��ev����Y;�uV���E����u�VW�f����V����_^[�Ë�V������W��;�s���t�Ѓ�;�r�_^Ë�V������W��;�s���t�Ѓ�;�r�_^Ë�U��QQV蚗�������F  �V\��W�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ���=����;�}$k��~\�d9 �=���B߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]Ë�U����\��e� �e� SW�N�@��  ��;�t��t	�У`��`V�E�P���u�3u�� �3��X�3����3��E�P����E�3E�3�;�u�O�@����u������5\��։5`�^_[�Ë�U���(3�S�]V�uW�}�E��E��E��E��E��E��E��E�9�t�5�}���Y���F�M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E�d���M��]�Q��]���]���Y����  �٘��� "   �  �E�`���M��]�Q��E�   �]���]���Y�j  �E�   �E�`���E�X���]���]���"  �M��E�X��r����E�T��׉M��E�T��Z����E�d�놃�tNIt?It0It ��t����   �E�L���E�D���E�d�����E�d��x����E�   ��������   �E�   �E�<���������������   �$�T��E�T���E�X���E�`���E�4���E�,���E�$��y����E���m����E����E����E����M����]���]�M��]�Q�E�   ��Y��u�A���� !   �E��_^[�û�����������s���]�T� �	���% 褙���3�Ë�U��QQSV���  V�5��gw  �EYY�M�ظ�  #�QQ�$f;�uU�v  YY��~-��~��u#�ESQQ�$j�t  ���rVS�w  �EYY�d�ES�x����\$�E�$jj�?�xu  �]��EY�]�Y����DzVS��v  �E�YY�"�� u��E�S���\$�E�$jj�pt  ��^[�Ë�U��E��]Ë�U���5�����Y��t�u��Y��t3�@]�3�]Ë�U��� S3�9]u �ȕ��SSSSS�    �H��������   �MV�u;�t!;�u處��SSSSS�    �H��������S�����E�;�w�M�W�u�E��u�E�B   �u�u�P�u��w  ����;�t�M�x�E����E�PS����YY��_^[�Ë�U���uj �u�u�u�5�����]�jhH��<���3��]3�;���;�u�����    WWWWW��G��������S�=|+u8j����Y�}�S�/���Y�E�;�t�s���	�u���u��E������%   9}�uSW�5�������������3��]�u�j�ԥ��Y������U���0���S�ٽ\�����=` t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=` t�#  ��8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����,  �   [�À�8�����=< uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ��������������x�����s4����,ǅr���   ��������������p�����v���VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�*�  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����D   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Àzuf��\���������?�f�?f��^���٭^������剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^������剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp��������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-���p��� ƅp���
��
�t����������l$�l$�D$���   5   �   t�������� u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t���������l$������������l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r ���������|$�l$�ɛ�l$������l$��Ã�,��?�$�>����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  ������� �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����,�Ƀ�u�\$0�|$(���l$�-4�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8��l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w����|$��<$� �|$$�D$$   �D$(�l$(����<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  ������� �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����,�Ƀ�u�\$0�|$(���l$�-4�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8��l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w����|$��<$� �|$$�D$$   �D$(�l$(����<$�l$$�Q�����0Z�����0Z�������@���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�p  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��̳������������������   s��ܳ��ĳ������������������   v��Գ떋�U����\�3ŉE�j�E�Ph  �u�E� ����u����
�E�P�D��Y�M�3��R*���Ë�U���4�\�3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5t��M�QP�֋l���t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u��$[����YF;�~[�����wS�D6=   w/������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�H��Y;�t	� ��  ���E���}�9}�t؍6PW�u��l)����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�h���t`�]��[�h�9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�[Y��YY�E�;�t+WWVPV�u�W�u��;�u�u��I2��Y�}���}��t�MЉ�u��t%��Y�E��e�_^[�M�3��(���Ë�U���S�u�M��j%���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P��8  YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP��  �� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U��QQ�\�3ŉE���SV3�W��;�u:�E�P3�FVh@�V����t�5��4�H���xu
jX���������   ;���   ����   �]�9]u��@�E�5l�3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�c}����;�t� ��  �P�)F��Y;�t	� ��  ���؅�ti�?Pj S��&����WS�u�uj�u�օ�t�uPS�u���E�S�y#���E�Y�u3�9]u��@�E9]u��@�E�u�����Y���u3��G;EtSS�MQ�uP�u��������;�t܉u�u�u�u�u�u����;�tV�/��Y�Ǎe�_^[�M�3��,&���Ë�U����u�M���"���u$�M��u �u�u�u�u�u�������}� t�M��ap���jhh������M3�;�v.j�X3���;E�@u�{���    WWWWW�.����3���   �M��u;�u3�F3ۉ]���wi�=|+uK������u�E;l+w7j詍��Y�}��u试��Y�E��E������_   �]�;�t�uWS�U%����;�uaVj�5��`���;�uL9=�t3V����Y���r����E;��P����    �E���3��uj�M���Y�;�u�E;�t�    ���K����jh��������]��u�u��C��Y��  �u��uS�.��Y�  �=|+��  3��}�����  j趌��Y�}�S�ߌ��Y�E�;���   ;5l+wIVSP���������t�]��5V萔��Y�E�;�t'�C�H;�r��PS�u��D��S菌���E�SP赌����9}�uH;�u3�F�u������uVW�5��`��E�;�t �C�H;�r��PS�u���C��S�u��h������E������.   �}� u1��uF������uVSj �5��������u�]j����YË}����   9=�t,V�_���Y��������Vy��9}�ul���H�P�y��Y��_����   �1y��9}�th�    �q��uFVSj �5��������uV9�t4V�����Y��t���v�V�����Y��x���    3��X������x���|�����u��x�����H�P�tx���Y���ҋ�U��MS3�;�v(j�3�X��;Es�x��SSSSS�    �{+����3��A�MVW��9]t�u�V���Y��V�u������YY��t;�s+�Vj �S�Y"������_^[]Ë�U��E��������]Ë�U��E��V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5���q��Y�j h������3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�~s�����}؅�u����a  �����`�w\���]���������Z�Ã�t<��t+Ht�Vw���    3�PPPPP�@*����뮾���������
�����E�   P�!q���E�Y3��}���   9E�uj����9E�tP�+���Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.���M܋����9M�}�M�k��W\�D�E����p����E������   ��u�wdS�U�Y��]�}؃}� tj 蹇��Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3�裓��Ë�U����HB�PD�M��U���u����Ãe� SW�E��FPj1Q3�C�E�SP��������FPj2�u��E�SP������FPj3�u��E�SP������FPj4�u��E�SP������P��FPj5�u��E�SP�u�����FPj6�u��E�SP�`���Vj7�u���E�SP�N�����F Pj*�u��E�SP�9�����P��F$Pj+�u��E�SP�!�����F(Pj,�u��E�SP������F,Pj-�u��E�SP�������F0Pj.�u��E�SP�������P��F4Pj/�u��E�SP�������FPj0�u��E�SP������F8PjD�u��E�SP������F<PjE�u��E�SP������P��F@PjF�u��E�SP�s�����FDPjG�u��E�SP�^�����FHPjH�u��E�SP�I�����FLPjI�u��E�SP�4�����P��FPPjJ�u��E�SP������FTPjK�u��E�SP������FXPjL�u��E�SP�������F\PjM�u��E�SP�������P��F`PjN�u��E�SP�������FdPjO�u��E�SP������FhPj8�u��E�SP������FlPj9�u��E�SP������P��FpPj:�u��E�SP�n�����FtPj;�u��E�SP�Y�����FxPj<�u��E�SP�D�����F|Pj=�u��E�SP�/�����P����   Pj>�u��E�SP��������   Pj?�u��E�SP���������   Pj@�u�S�E�P���������   PjA�u��E�SP�������P����   PjB�u��E�SP��������   PjC�u��E�SP��������   Pj(�u��E�SP��������   Pj)�u��E�SP�i�����P����   Pj�u��E�SP�N�������   Pj �u��E�SP�6�������   Ph  �u��E�SP��������   Ph	  �]�S�E�j P�������P���_���   [�Ë�U��V�u����  �v�l%���v�d%���v�\%���v�T%���v�L%���v�D%���6�=%���v �5%���v$�-%���v(�%%���v,�%���v0�%���v4�%���v�%���v8��$���v<��$����@�v@��$���vD��$���vH��$���vL��$���vP��$���vT��$���vX�$���v\�$���v`�$���vd�$���vh�$���vl�$���vp�$���vt�$���vx�z$���v|�r$����@���   �d$�����   �Y$�����   �N$�����   �C$�����   �8$�����   �-$�����   �"$�����   �$�����   �$�����   �$�����   ��#����,^]Ë�U��SVW�}�  �@t@h�   j�J����YY��u3�@�E��������tV�+���V�#��YY��ǆ�      �����   �;�t�   P���73�_^[]Ë�U��V�u��t5�; tP�Z#��Y�F;tP�H#��Y�v;5tV�6#��Y^]Ë�U���S�]V3�W�]�u�9su9su�u��u��E �:  j0j��I����YY�};�u3�@�w  ���   jYj��|I��3�Y�E�;�u�u��"��Y�щ09s��   j�UI��Y�E�;�u3�F�u�"���u��"��YY���  �0�u�{>VjW�E�jP������E�FPjW�E�jP�����	E�FPjW�E��E�jP������<E�tV����Y���뎋E�� ����0|��9��0�@�8 u��7��;u���~�����> u��� �E���H��u��H�E�3�A��E���t����   �5���tP�֋��   ��tP�օ�u���   �!�����   �!��YY�E����   �E����   �E���   3�_^[�Ë�U��V�u��t~�F;tP�J!��Y�F;tP�8!��Y�F;tP�&!��Y�F;tP�!��Y�F;tP�!��Y�F ; tP�� ��Y�v$;5$tV�� ��Y^]Ë�U���SV�uW3��}��u��}�9~u9~u�}��}�� �6  j0j�G����YY;�u3�@�u  j�1G��Y�E�;�u	S�y ��Y���89~��  j�G��Y�E�;�uS�V ���u��N ��Y�҉8�v8�CPjV�E�jP�������CPjV�E�jP������CPjV�E�jP�s�����CPjV�E�jP�_�����P��CPjV�E�jP�H�����C PjPV�E�jP�4�����C$PjQV�E�jP� �����C(PjV�E�j P������P��C)PjVj �E�P�������C*PjTV�E�j P�������C+PjUV�E�j P�������C,PjVV�E�j P������P��C-PjWV�E�j P������C.PjRV�E�j P������C/PjSV�E�j P�z�����<�t$S����S�����u������u��������Q����C����0|��9��0�@�8 u��#��;u���~�����> u���jY� ���E�u�   ��	���I�K� �@�M��C3�@3��9}�t�M�����   ;�tP�����   ;�t#P����u���   �@�����   �5��YY�E����   �E����   ���   3�_^[�Ë�U��ES3�VW;�t�};�w�yj��j^�0SSSSS�f�������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u��2j��j"Y����3�_^[]��������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^�Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w�i��j^�0SSSSS���������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x�����#i��j"Y���낋�U��3�S3�@9]|FVW��t>�EÙ+��E���<��7�E�0��X  YY��u
�M���9�}N�u��^;]~�_^3Ʌ���[��]Ë�U����\�3ŉE�V���tS�> tNh��V�Z��YY��t=h�V�Z��YY��uj�E�Pj�w����t/�u�V�,��Y�M�3�^�N����j�E�Ph  �w����u3��׍E�h�P�MZ��YY��u��x�뻋�U��3�f�Mf;�ؼt@@��r�3�@]�3�]Ë�V3��#��,aB<w������,A<w��������tЊ
��u׋�^�3��
B��A|��Z~��a��w@��Ë�U���|�\�3ŉE�VW�}��c�����ׁƜ   ������jx�E�P�F���%���  PW����u!F@�2�E�P�v�UW  YY��uW����Y��t
�N�~�~�F���Ѓ��M�_3�^����� ��U���|�\�3ŉE�Vjx�E�P�E%�  j   P������u3��.�U������9Et�} t�6W�������V���B��Y;�_t�3�@�M�3�^����Ë�U���|�\�3ŉE�SVW�}��b�����ׁƜ   �y�������jx�E�P�F���%���  PW�Ӆ�u�f 3�@�b  �E�P�v�@V  YY����   jx�E�P�F���%���  PW�Ӆ�t��E�P�6�V  YY��u�N  �~�R�FuO�F��t,P�E�P�6�%W  ����u�6�N�~�A��Y;Fu!�~��V��uW����Y��t	���V�~�N�   #�;���   jx�E�P�F���%���  PW�Ӆ������E�P�6�eU  Y3�Y��u/�N   �F9^t
   �F�G9^t;�6�}@��Y;Fu.j�9^u49^t/�E�P�6�U  YY��uSW�������YY��t�N   9^u�~�F���Ѓ��M�_^3�[������ ��U���|�\�3ŉE�VW�}�a�����ׁƜ   ������jx�E�P�F���%���  PW����u!F@�[�E�P�6�xT  YY��u	9Fu0j��~ u0�~ t*�E�P�6�RT  YY��uPW���$���YY��t
�N�~�~�F���Ѓ��M�_3�^����� �6�V?���v�����@�F�C?��������f @�~ YY�FtjX���	���jh���F���F�   t�   t�u�f ��6��>�������@Y�FtjX������jh� �F���Fu�f Ë�U��SVW�_���]���Ɯ   ��u�N  �   �C@�~����t�8 tWjh ����������f ��tS�8 tN���t�8 t�������S����~ ��   Vj@h���������tb�?��t�? t�����P�����I�?��t0�? t+W�>������Y�j@h���F���Fu�f ��F  ���F�F�~ ��   �˃����#ˋ��������}����   ����  ��   ����  ��   ��P�������   j�v� �����   �E��tf�Nf�f�Nf�Hf�x�]��tm�=��  f9u%h��j@S�b������t"3�PPPPP������j@Sh  �v�ׅ�t,j@�C@Ph  �v�ׅ�tj
j��S�u�T  ��3�@�3�_^[]Ë�U��VW�}�ǃ� ��  H��  H��  H�I  H��  �M�ESj Z�r  �0;1t|�0�+�t3ۅ��Í\�����i  �p�Y+�t3ۅ��Í\�����H  �p�Y+�t3ۅ��Í\�����'  �p�Y+�t3ۅ��Í\����3����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3����r  �p;qt~�p�Y+�t3ۅ��Í\�����I  �p	�Y	+�t3ۅ��Í\�����(  �p
�Y
+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����w  �p�Y+�t3ۅ��Í\����3����R  �p;qt~�Y�p+�t3ۅ��Í\�����)  �p�Y+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����x  �p�Y+�t3ۅ��Í\�����W  �p�Y+�t3ۅ��Í\����3����2  �p;qt~�p�Y+�t3ۅ��Í\�����	  �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\����3�����   �p;qtr�p�Y+�t3ۅ��Í\����u}�p�Y+�t3ۅ��Í\����u`�p�Y+�t3ۅ��Í\����uC�p�Y+�t3ۅ��Í\����3���u"��+�;�������σ���  �$�����  �P�;Q�tq���Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����3����v����P�;Q�t}���Q�+�t3҅��T�����N����p��Q�+�t3҅��T�����-����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����}����p��Q�+�t3҅��T����3����X����P�;Q�t}���Q�+�t3҅��T�����0����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T�����^����p��Q�+�t3҅��T����3����9����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�to���Q�+�t3҅��T���u6�p��Q�+�t3҅��T���u�p��Q�+�t3҅��T���t����@��I�+�t3Ʌ����L	����3���u3�[�S  �P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����n����p��Q�+�t3҅��T�����M����p��Q�+�t3҅��T�����,����p��Q�+�t3҅��T����3��������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����x����P�;Q�t}���Q�+�t3҅��T�����P����p��Q�+�t3҅��T�����/����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3����Z����P�;Q�t~�Q��p�+�t3҅��T�����1����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����`����p��Q�+�t3҅��T����3����;����I��@�+�� ���3Ʌ����L	���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����b����p��Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����l����P�;Q�t}���Q�+�t3҅��T�����D����p��Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����s����p��Q�+�t3҅��T����3����N����P�;Q�t~�Q��p�+�t3҅��T�����%����Q��p�+�t3҅��T���������Q��p�+�t3҅��T����������Q��p�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T����3����/���f�P�f;Q�������Q��p�+������3҅��T����  �����P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����i����P�;Q�t}���Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����p����p��Q�+�t3҅��T����3����K����P�;Q�t}���Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T�����r����p��Q�+�t3҅��T�����Q����p��Q�+�t3҅��T����3����,����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T�����3����p��Q�+�t3҅��T����3��������p��Q�+������3҅��T���������������M�u��+�t3҅��T�����   �A�V+�t3҅��T�����   �A�V+�t3҅��T�����   �A�N+���   3Ʌ����L	����   �M�u��+�t3҅��T���uh�A�V+�t3҅��T���uK�A�N랋M�u��+�t3҅��T���u �A�N�p����E�M� �	�_���3�_^]ø���;'H�����)�
my��	��o	O[|�������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U�����SV�uW3��E��}�}��}��FFf�> t����at8��rt+��wt�cJ��WWWWW�    �O�����3��S  �  �3ۃM��	�	  �M�3�AFF�f;���  � @  ;��   ����S��   ��   �� ��   ��tVHtG��t1��
t!���u���9}���   �E�   ����   �ˀ   �   ��@��   ��@�   �E�   �   ����   �E����������   �E��}9}�ur�E�   �� �l��TtX��tCHt/��t��������� �  uC��E9}�u:�e������E�   �09}�u%	U��E�   ��� �  u�� �  ��   ��t3���FF�f;������9}���   �FFf�> t�jVh��.E  �����`���j ��X�FFf9t�f�>=�G���FFf9t�jh�V�PD  ����u��
��   �Djh �V�1D  ����u����   �%jh4�V�D  �������������   �FFf�> t�f9>�����h�  �u�ES�uP��B  ����������E�@�M��H�M�x�8�x�x�H_^[��jh��� e��3�3��}�j�Z��Y�]�3��u�;5`+��   �@��9t[� �@��uH� �  uA�F���w�FP�Y��Y����   �@�4�V�]u��YY�@���@�tPV�u��YYF둋��}��h��j8�y!��Y�@��@�9tIh�  � �� P�  YY���@u�4����Y�@����� P�(��@�<�}�_;�t�g �  �_�_��_�O��E������   ���Fd��Ë}�j�#X��Y�SVW�T$�D$�L$URPQQh\d�5    �\�3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�
  �   �C�
  �d�    ��_^[ËL$�A   �   t3�D$�H3��	���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j��	  3�3�3�3�3���U��SVWj j h Q�i  _^[]�U�l$RQ�t$������]� ��U����u�M��5����E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]�������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �������U��W�}3�������ك��E���8t3�����_�Ë�U���SV�u�M������]�   ;�sT�M胹�   ~�E�PjS������M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P����YY��t�Ej�E��]��E� Y��D��� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�����$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=d u�E�H���w�� ]�j �u�����YY]Ë�U���(�\�3ŉE�SV�uW�u�}�M��3����E�P3�SSSSW�E�P�E�P��J  �E�E�VP�H@  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[������Ë�U���(�\�3ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P�5J  �E�E�VP��D  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�)����Ë�U��MSV�u3�W�y;�u�B��j^�0SSSSS����������   9]v݋U;ӈ~���3�@9Ew��A��j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W����@PWV������3�_^[]Ë�U��Q�M�ASVW������  #�% �  �߉E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��E��<  �U����������U��E�����P������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0�\�3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��O  �uЉC�E։�EԉC�E�P�uV�������$��t3�PPPPP�������M�_�s^��3�[�"����������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j賛��YË�U��E�M%����#�V������t1W�}3�;�tVV��W  YY���>��j_VVVVV�8���������_��uP�u��t	�W  ���W  YY3�^]Ë�U��E�]�jh����[���e� �u�u�$��E��/�E� � �E�3�=  �����Ëe�}�  �uj����e� �E������E��[���������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h�h �d�    P��SVW�\�1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U��3�@�} u3�]��U��SVWUj j h�(�u�`  ]_^[��]ËL$�A   �   t2�D$�H�3�����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�(d�5    �\�3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�(u�Q�R9Qu�   �SQ�@�SQ�@�L$�K�C�kUQPXY]Y[� ���jh(��X��3ۉ]�j�M��Y�]�j_�}�;=`+}W�����@�9tD� �@�tP����Y���t�E��|(�@��� P�$��@�4����Y�@�G��E������	   �E��yX���j�YL��YË�U����UV�uj�X�E�U�;�u��:���  ��:��� 	   ����  S3�;�|;5 r'�:����:��SSSSS� 	   ����������Q  ����W�<�@�����ƊH��u�q:����W:��� 	   �j�����wP�]�;��  ����  9]t7�@$����E���HjYtHu���Шt����U�E�E��   ���Шu!�:�����9���    SSSSS��������4����M;�r�E�u����Y�E�;�u�9���    �9���    ����h  jSS�u�^  ��D(�E���T,���AHtt�I��
tl9]tg��@�M�E�   �D
8]�tN��L%��
tC9]t>��@�M�}��E�   �D%
u$��L&��
t9]t��@�M�E�   �D&
S�M�Q�uP��4�ؐ���{  �M�;��p  ;M�g  �M��D� ���  �}��  ;�t�M�9
u��� ��]�E�É]�E�;���   �M�<��   <t�CA�M�   �E�H;�s�A�8
u
AA�M�
�u�E�m�Ej �E�Pj�E�P��4�ؐ��u
�H���uE�}� t?��DHt�}�
t����M��L�%;]�u�}�
t�jj�j��u�  ���}�
t�C�E�9E�G������D� @u����C��+E�}��E���   ����   K���xC�   3�@�����;]�rK�@��P t�����P��u�^7��� *   �zA;�u��@���AHt$C���Q|	���T%C��u	���T&C+���ؙjRP�u��  ���E�+]���P�uS�u�j h��  �l��E���u4�H�P�7��Y�M���E�;EtP�H���Y�E�����  �E��  �E��3�;�����E��L0��;�t�M�f�9
u��� ��]�E�É]�E�;���   �E�f����   f��tf�CC@@�E�   �M����;�s�Hf�9
u���Ej
�   �M�   �Ej �E�Pj�E�P��4�ؐ��u
�H���u[�}� tU��DHt(f�}�
t�jXf���M��L��M��L%��D&
�*;]�uf�}�
t�jj�j��u�|  ��f�}�
tjXf�CC�E�9E�������t�@u��f� f�CC+]�]������H�j^;�u�W5��� 	   �_5���0�i�����m�Y����]��\���3�_[^��jhH��\R���E���u�'5���  �5��� 	   ����   3�;�|; r!��4���0��4��� 	   VVVVV��������ɋ�����@��������L9��t�����;M�Au�4���0�4���    �P��  Y�u���D8t�u�u�u�~������E���`4��� 	   �h4���0�M���E������	   �E��Q����u�  YË�U��QQ�EV�u�E��EWV�E���  ���Y;�u�4��� 	   �ǋ��J�u�M�Q�u�P�ܐ�E�;�u�H���t	P��3��Y�ϋ�����@�����D0� ��E��U�_^��jhh���P������u܉u��E���u�3���  �3��� 	   �Ƌ���   3�;�|; r!�r3���8�X3��� 	   WWWWW�D������ȋ�����@��������L1��u&�13���8�3��� 	   WWWWW������������[P�=  Y�}���D0t�u�u�u�u�������E܉U����2��� 	   ��2���8�M���M���E������   �E܋U��P����u�z  YË�U��E���u�2��� 	   3�]�V3�;�|; r�b2��VVVVV� 	   �N�����3���ȃ�����@���D��@^]Ë�U����\�3ŉE�V3�95PtO�=�
�u�N  ��
���u���  �pV�M�Qj�MQP�0���ug�=Pu��H���xuω5PVVj�E�Pj�EPV�,�P�h���
���t�V�U�RP�E�PQ�(���t�f�E�M�3�^�w������P   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M������E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�l����E�u�M;��   r 8^t���   8]��e����M��ap��Y����0��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�l����:���뺋�U��j �u�u�u�������]Ë�U��EVW��|Y; sQ���������<�@����<�u5�=XS�]u�� tHtHuSj��Sj��Sj��4���3�[���/��� 	   ��/���  ���_^]Ë�U��MS3�;�VW|[; sS������<�@�������@t5�8�t0�=Xu+�tItIuSj��Sj��Sj��4����3���F/��� 	   �N/������_^[]Ë�U��E���u�2/���  �/��� 	   ���]�V3�;�|"; s�ȃ�����@����@u$��.���0��.��VVVVV� 	   ������������ ^]�jh����K���}����������4�@�E�   3�9^u6j
��@��Y�]�9^uh�  �FP�����YY��u�]��F�E������0   9]�t����������@�D8P�(��E��K���3ۋ}j
�?��YË�U��E�ȃ�����@���DP�,�]�jh���"K���M��3��}�j�V?��Y��u����b  j�@��Y�}��}؃�@�<  �4�@����   �u���@   ;���   �Fu\�~ u9j
�?��Y3�C�]��~ uh�  �FP�����YY��u�]���F�e� �(   �}� u�^S�(��FtS�,���@낋}؋u�j
�>��YÃ}� u��F��+4�@��������u�}��uyG�+���j@j �N��YY�E���ta��@��  ���   ;�s�@ ���@
�` ��@�E������}�����σ�����@�DW�����Y��u�M���E������	   �E���I���j��=��Y�����V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U���SVW�%���e� �= ����   h���8������*  �5��h��W�օ��  P�%���$��W���P��$���$��W���P��$���$h�W� ��P��$��Y�(��thP�W��P�$��Y�$�$;�tO9(tGP�	%���5(����$��YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9�;�t0P�$��Y��t%�ЉE���t� ;�tP�$��Y��t�u��ЉE��5�$��Y��t�u�u�u�u����3�_^[�Ë�U��MV3�;�|��~��u�T�(�T�T��%*��VVVVV�    ���������^]Ë�U����u�M�������u�u�u�u�<��}� t�M��ap��Ë�U��QQ�\�3ŉE��,S�<�VW3�3�G;�u,VVWV�Ӆ�t�=,�/�H���xu
jX�,��,����   ;���   ;�u#9uu�E� �@�EVV�u�u�ӋȉM�;�u3��   ~Ej�3�X���r9�D	=   w�r)����;�t����  ���P�5���Y;�t	� ��  �����3�;�t��u�W�u�u�Ӆ�t VV9uuVV��u�uj�WV�u�h���W����Y����u�u�u�u���e�_^[�M�3������Ë�U����u�M��h����u�E��u�u�u�uP�������}� t�M��ap��Ë�U��E�0]Ë�U����u�M������E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u�D��M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�}  Y����  �t�Etj�c  Y����v  ����   �E��   j�A  �EY�   #�tT=   t7=   t;�ub��M����`	��{L�H��M�����{,�`	�2��M�����z�`	���M�����z�P	��P	��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�x  �M��]�� �����������}�E���P��S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}��"��� "   ]���"��� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���h;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�s������uV�,���Y�E�^�Ë�l�h��  �u(�  �u�����E ���Ë�U��=` u(�u�E���\$���\$�E�$�uj�/�����$]���!��h��  �u� !   �J  �EYY]Ë�S��QQ�����U�k�l$���   �\�3ŉE��s �CP�s��������u"�e���CP�CP�s�C �sP�E�P�I������s�p������=` u+��t'�s �C���\$���\$�C�$�sP�r�����$�P�����$��  �s �  �CYY�M�3��������]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj���  f;�u�E�� u9Utj��3�]Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������"Q���EQQ�$����������  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�-x	�]���t����-x	�]�������t
�-�	�]����t	�������؛�� t���]����jh���<��3�9�+tV�E@tH9�	t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�	 �e��U�E�������e��U��;����A@t�y t$�Ix��������QP��P��YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u�����8*u�ϰ?�d����} �^[]Ë�U���x  �\�3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������J�����u5�_���    3�PPPPP�I����������� t
�������`p������
  �F@u^V�lO��Y�����t���t�ȃ��������@����A$u����t���t�ȃ������@����@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw����0���3��3�3����P�j��Y������;���	  �$�.S��������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�����������Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u��	������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P�d6  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  ��	������P�_���Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7����������3  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V� ���������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5�����Y�Ћ���������   t 9�����u������PS�5���c��Y��YY������gu;�u������PS�5���>��Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�q�����0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u��	�������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF��0  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t�������+��������� Y���������������t������������������������� t
�������`p��������M�_^3�[�Z����Ð9K:IjI�IJJeJ�K��S��QQ�����U�k�l$���   �\�3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|�����������uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�;�����h��  ��x���������>YYt�=` uV�Q���Y��u�6����Y�M�_3�^�������]��[Ë�U��UV�uW��H�F��w�� �
�y�B��w�� ��t;�t�_+�^]Ë�U���S�u�M�荷��3�9]u.���SSSSS�    ������8]�t�E��`p������   W�};�u+�i��SSSSS�    �U�����8]�t�E��`p������U�E�9XuW�u�:���YY�4V�E� �M�QP�e����E����M�QP�S�����G;�t;�t�+���^8]�t�M��ap�_[�Ë�U��V3�95du09uu����VVVVV�    �����������9ut�^]����V�u�u�������^]Ë�U���S3�VW9]��   �u�M��Y���9]u.�m��SSSSS�    �Y�����8]�t�E��`p������   �};�t˾���9uv(�.��SSSSS�    ������8]�t�E��`p����`�E�9Xu�uW�u��,  ��8]�tD�M��ap��;�E� �M�QP�����E����M�QP������G�Mt;�t;�t�+����3�_^[�Ë�U��V3�95du99uu���VVVVV�    �x����������'9ut܁}���w�^]�H,  V�u�u�u������^]Ë�U��QSV��3�;�u�3��j^SSSSS�0� ��������   W9]w���j^SSSSS�0����������   3�9]���A9Mw	����j"�ЋM�����"w��]���9]t�-�N�E�   �؋�3��u��	v��W���0�A�E�3�;�v�U9U�rڋE�;Er�럈I���I�G;�r�3�_^[�� ��U��}
�Eu
��}jj
�j �u�u�M�����]Ë�U���4S3��E�VW���]��]��E�   �]�t	�]��E��
�E�   �]��E�P�-  Y��tSSSSS�ž�����M� �  ��u�� @ u9E�t�M������+ú   ��   �tGHt.Ht&����������j^SSSSS�0薿�����  �U����t��   u��E�   @��}��EjY+�t7+�t*+�t+�t��@u�9}����E���E�   ��E�   ��E�   ��]��E�   #¹   ;��   ;t0;�t,;�t=   ��   =   �@����E�   �/�E�   �&�E�   �=   t=   t`;������E�   �E�E�   ��t�h��#M��x�E�   �@t�M�   �M�   �M��   t	}�� t�M�   ��E�   릨t�M�   �c�������u�]������@���    �   �E�=@�S�u��    �u�E�P�u��u��u�׉E���um�M��   �#�;�u+�Et%�e����S�u�E��u�P�u��u��u�׉E���u4�6������@�����D0� ��H�P��
��Y�
��� �u  �u����;�uD�6������@�����D0� ��H���V�
��Y�u�� �;�u��R
���    룃�u�M�@�	��u�M��u��6�������Ѓ�����@Y��Y�M����L��Ѓ�����@���D$� ��M��e�H�M���   �����  �Etrj���W�6�J�����E�;�u��	���8�   tN�6�_N�������j�E�P�6�]���������uf�}�u�E�RP�6��'  ��;�t�SS�6�FJ����;�t��E���0  � @ � @  �}u�E�#�u	M�	E�E#�;�tD=   t)= @ t"=   t)= @ t"=   t= @ u�E���M�  #�;�u	�E���]��E   ��  �E�@�]���  �E��   �#�=   @��   =   �tw;���  �E�;��y  ��v��v0���f  �E�3�H�&  H�R  �E���  �E�   �  jSS�6�*������t�SSS�6����#���������j�E�P�6�?���������t�����tk����   �}�﻿ uY�E���   �E�;���   ���b������P���jSS�6��������C���SSS�6������#����   �����E�%��  =��  u�6�TL��Y���j^�0���d  =��  uSj�6�XH�������������E��ASS�6�=H������E�﻿ �E�   �E�+�P�D=�P�6�B������������9}�ۋ������@�����D$�2M���0�������@�����D$�M�������
ʈ8]�u!�Et��ȃ�����@���D� �}��   ���#�;�u|�Etv�u�� �S�u�E�jP�u������W�u�@����u4�H�P�����ȃ�����@���D� ��6����Y�����6������@�������_^[��jh���P#��3��u�3��};���;�u����j_�8VVVVV���������Y��3�9u��;�t�9ut�E%������@tu��u�u�u�u�E�P���i������E��E������   �E�;�t���	#���3��}9u�t(9u�t�����������@�D� ��7�=���YË�U��j�u�u�u�u�u������]Ë�U���SV3�3�W9u��   �];�u"���VVVVV�    ������������   �};�t��u�M��ī���E�9pu?�f��Ar	f��Zw�� ���f��Ar	f��Zw�� CCGG�M��tBf��t=f;�t��6�E�P�P�%  ���E�P�P�u%  ��CCGG�M��t
f��tf;�t�����+��}� t�M��ap�_^[�Ë�U��V3�W95du3�9u��   �};�u�#��VVVVV�    �����������`�U;�t��f��Ar	f��Zw�� ���f��Ar	f��Zw�� GGBB�M��t
f;�tf;�t�����+��V�u�u�u�w�����_^]Ë�U��} u3�]ËU�M�Mt�f��tf;uAABB����
+�]Ë�U����  ��f9Eu�e� �e�   f9Es�E���f�Af#E���E��@�u�M������E��p�p�E�Pj�EP�E�jP�$  ����u!E��}� t�E�`p��E��M#��Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5X
N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�T
��+X
;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5X
N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��\
A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;P
�\
��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�P
�d
�3�@�   �d
�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+\
��M���Ɂ�   �ً`
]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5p
N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�l
��+p
;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5p
N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��t
A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;h
�t
��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�h
�|
�3�@�   �|
�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+t
��M���Ɂ�   �ًx
]���@u�M�U�Y��
�� u�M�_[�Ë�U���|�\�3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u����SSSSS�    �������3��O  �U�U��< t<	t<
t<uB��0�B���/  �$��s�Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �#  =�����/  ��
��`�E�;���  }�عP�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9U�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �;����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[薛�����mnmn�n�no1o�owo�o�o�o��U���t�\�3ŉE�S�]VW�u�}�f��E��U�� �  #��E��A�#�f�}� �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   t�C-��C �u�}�f��u1��u-��u)3�f9M�f�����$ �C�C�C0�C 3�@�  f;���   3�@f��   �;�u��t��   @uh��Sf�}� t��   �u��u;h���;�u0��u,h���CjP������3���tVVVVV�
������C�*h���CjP赙����3���tVVVVV�ޡ�����C3��s  �ʋ�i�M  �������Ck�M��������3���f�M��
�ۃ�`�E�f�U�u�}�M�����  }�P�ۃ�`�E�����  �E�T�˃������h  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��z����M�����?  ��  f;���  �]��E�3��ɉU��U��U�U��U�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��U���3�3�f9u���H%   � ���E��[���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �_�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[�|����À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95�+��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E������Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��3�PPjPjh   @h��D���
á�
V�5 ����t���tP�֡�
���t���tP��^á\���3�9�����Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v�\���j^SSSSS�0�I��������V�u�M������E�9X��   f�E��   f;�v6;�t;�vWSV�,������	���� *   ������ 8]�t�M��ap�_^[��;�t2;�w,�����j"^SSSSS�0�˕����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�h�;�t9]�^����M;�t����H���z�D���;��g���;��_���WSV�U������O�����U��j �u�u�u�u�|�����]�U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U���SVW3�jSS�u�]��]��e����E�#��U���tYjSS�u�I�����#ʃ����tA�u�}+����   ;���   �   Sj�L�P�`��E���u�2����    �'���� _^[��h �  �u�  YY�E���|
;�r�����P�u��u��������t6�+��xӅ�wϋu��u��u��   YY�u�j �L�P�L�3��   ������8u�����    ����u��;�q|;�skS�u�u�u�N���#�����D����u�7���YP�H������H��E�#U���u)�F����    �N������H���u�#u��������S�u��u��u����#���������3��������U��S�]V�u������@������0�A$�W�y����   ���� @  tP�� �  tB��   t&��   t��   u=�I��
�L1$��⁀���'�I��
�L1$��₀���a��I��
�L1$�!���_^[u� �  ]����% �   @  ]Ë�U��EV3�;�u�.���VVVVV�    ������jX�
� �3�^]Ë�U����  �ȃ�f9M��   S�u�M��ƅ���M�Q3�;�u�E�H�f��w�� ���aV�   ��f9u^s)�E�Pj�u�9��������Et9�M싉�   f����q�M�jQj�MQPR�E�P�*  �� ���Et�E�8]�t�M�ap�[�Ë�U����u�M��#����}�}3���u�u�u�u���}� t�M��ap��Ë�U����\�3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[�J����Ë�U����u�M������E��~�M��Jf�9 t	AA��u���+�H�u �uP�u�u�u�p��}� t�M��ap����%P������̋T$�B�J�3��ԅ���p��c�������̋T$�B�J�3�贅������C�������̋T$�B�J�3�蔅���T��#�������̋T$�B�J�3��t��������������̋T$�B�J�3��T�������������̋T$�B�J�3��4�������Ï������̋T$�B��h���3������J�3��������閏���������̋T$�B�����3������4��p����̋T$�B�J�3��Ą������S�������̋T$�B�J�3�褄���@��3�������̋T$�B�J�3�脄���J�3��z�������	�������������̋T$�B�J�3��T��������������̋T$�B�J�3��4����H��Î������̋T$�B�J�3��������风������̋T$�B�J�3������J�3��������y�������������̋T$�B�J�3��ă������S�������̋T$�B�J�3�褃������3�������̋T$�B�J�3�脃���@������M��]w���T$�B�J�3��a������������M�����T$�B�J�3��>�������͍���M�����M��������T$�B�J�3��������韍���M���v���u��n��YËT$�B�J�3������(��r����M�鼇���T$�B�J�3�������T��O����T$�B�J�3�襂���@��4���������h@�����Yù���u��h�������Y�h������Yù8��u��h���ڦ��Y�h���Φ��YÃ=� uK����t���Q<P�B�Ѓ���    ����tV�������V�
m������    ^ù��u�����G���8�lu���9�}��                                                                   �� �� �� �� �� ,� D� \� d� �� �� �� �� �� �� � *� >� P� `� l� x� �� �� �� �� �� �� �� � � � (� :� N� `� n� z� �� �� �� �� �� �� �� �� �� �  � .� @� L� \� n� �� �� �� �� �� �� �� � *� D� T� j� �� �� �� �� �� �� �� � *� :� P� `� p� �� �� �� �� ��     �         ���4����        �3�^�hR���        ���                    {qP       �   �� �� bad allocation  @�P" � �  ��  �    0�3D-COAT     c:\program files\maxon\cinema 4d r13\plugins\applink_cinema4d\source\applinkdialog.cpp  Start import!   To import a new object? File exists!    export.txt  Folder ..\MyDocuments\3D-CoatV3\Exchange not found! 3D-CoatV3   Exchange    preference.ini  3D-Coat.exe is run! 3D-Coat.exe not found!  open    Start export!               c:\program files\maxon\cinema 4d r13\plugins\applink_cinema4d\source\applinkexporter.cpp    
   c:\program files\maxon\cinema 4d r13\resource\_api\ge_dynamicarray.h    ]   autopo  curv    prim    alpha   vox retopo  ref uv  ptex    mv  ppp [   # end   v       # begin      vertices
            �?vt   texture vertices
  /   f   usemtl   faces
 g   mtllib  mtl map_    illum 2
    Tr 0.000000
    Ns 50.000000
   Ks  Kd  Ka 0.300000 0.300000 0.300000
  newmtl  No selected objects!    Object "    " has no UVW tag.
UV coordinates can't be exported. Material not found on   object. Default Name    Export object   #Cinema4D Version:  %d.%m.%Y  %H:%M:%S  #File created:  #Wavefront OBJ Export for 3D-Coat
  File     write success! [SkipExport]
   [SkipImport]
         �import.txt  output.obj  obj ���� @�@� ��p� �� x�p� ����  �  � p� P� �� �� �� 0�  � `�       Y@��@�� ��  � � ��  � @
�
�� �� @�  � P� $���  � ` ��  � @
�
�  @�  � P� p�@� p� �� �� PPp�Selection   Error on inserting phongTag. Object:    Poly count:     V count:    Create objects...   Memory allocation error for material.   ����3@&� � P � @
�
�)�*`pp?d�����0�����L�0�vector<T> too long  bad cast    ios_base::eofbit set    ios_base::failbit set   ios_base::badbit set    ���E    X       P    can not removed!   normalmap   displacement %f displacement    map_Ks %s   map_Ks  map_Kd %s   map_Kd  Ke %lf %lf %lf  Ke  Ks %lf %lf %lf  Ks  Ka %lf %lf %lf  Ka  Kd %lf %lf %lf  Kd  illum %d    illum   d %lf   d   Ns %lf  Ns  newmtl %s   Open file   .    not found! c:\program files\maxon\cinema 4d r13\plugins\applink_cinema4d\source\applinkimporter.cpp    Nb faces:   Nb Grp:     Wrong face in OBJ file! f   vt  Gathering of data...        �dy���=vt %lf %lf %lf  vt %lf %lf  v %lf %lf %lf   g %s    mtllib %s   Parse file...   Open file:  textures.txt    `��W�V0�@��P��� �icon_coat.tif       c:\program files\maxon\cinema 4d r13\plugins\applink_cinema4d\source\applinkpreferences.cpp ���)�)�)�)�)�)�W          �?���^0j k�d`p`�ec:\program files\maxon\cinema 4d r13\resource\_api\c4d_file.cpp      �f@-DT�!	@D�0�п� �� �0��0��������������     @�@X�0�п� �� �0��0���������P�`��� �p�@���`�c:\program files\maxon\cinema 4d r13\resource\_api\c4d_gui.cpp  ��0�п� �� �0��p�8�0�п� �� �0��P����������� ����`�p� �P�Progress Thread 0%  ~   %       c:\program files\maxon\cinema 4d r13\resource\_api\c4d_general.h    %s         ����MbP?��P��r�0�    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_baseobject.cpp   c:\program files\maxon\cinema 4d r13\resource\_api\c4d_resource.cpp #   M_EDITOR    P���res c:\program files\maxon\cinema 4d r13\resource\_api\c4d_pmain.cpp        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_basetime.cpp      �Ngm��C   ����A  4&�k�  4&�kCd��� � �)�)    c:\program files\maxon\cinema 4d r13\resource\_api\c4d_libs\lib_ngon.cpp        c:\program files\maxon\cinema 4d r13\resource\_api\c4d_basebitmap.cpp   ��� c:\program files\maxon\cinema 4d r13\resource\_api\c4d_gv\ge_mtools.cpp �� <�� ��`���*   C   �����	�string too long invalid string position r            
   !   "   2   *            #   3   +       w   a   r b     w b     a b     r +     w +     a +     r + b   w + b   a + b   l�{��nUnknown exception   ���csm�               �                      �?      �?3      3            �      0C       �       ��                                                                                                                                                                                                                                                                                                        ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������LC_TIME LC_NUMERIC  LC_MONETARY LC_CTYPE    LC_COLLATE  LC_ALL  ��    �F|�8��Fp�8��;d�8�)�X�8���P�8��	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ _., _   ;   =   =;  EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    �e+000          �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    ʆ�Մbad exception   runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:    CorExitProcess  m s c o r e e . d l l         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow         �������             ��      �@      �              �?5�h!���>@�������             ��      �@      �        HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun united-states   united-kingdom  trinidad & tobago   south-korea south-africa    south korea south africa    slovak  puerto-rico pr-china    pr china    nz  new-zealand hong-kong   holland great britain   england czech   china   britain america usa us  uk  swiss   swedish-finland spanish-venezuela   spanish-uruguay spanish-puerto rico spanish-peru    spanish-paraguay    spanish-panama  spanish-nicaragua   spanish-modern  spanish-mexican spanish-honduras    spanish-guatemala   spanish-el salvador spanish-ecuador spanish-dominican republic  spanish-costa rica  spanish-colombia    spanish-chile   spanish-bolivia spanish-argentina   portuguese-brazilian    norwegian-nynorsk   norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg   german-lichtenstein german-austrian french-swiss    french-luxembourg   french-canadian french-belgian  english-usa english-us  english-uk  english-trinidad y tobago   english-south africa    english-nz  english-jamaica english-ire english-caribbean   english-can english-belize  english-aus english-american    dutch-belgian   chinese-traditional chinese-singapore   chinese-simplified  chinese-hongkong    chinese chi chh canadian    belgian australian  american-english    american english    american    �ENU ��ENU �ENU عENA йNLB ĹENC ��ZHH ��ZHI ��CHS ��ZHH ��CHS x�ZHI d�CHT T�NLB @�ENU 4�ENA $�ENL �ENC �ENB ��ENI �ENJ ܸENZ ĸENS ��ENT ��ENG ��ENU ��ENU t�FRB d�FRC P�FRL @�FRS 0�DEA �DEC �DEL ��DES �ENI طITS ̷NOR ��NOR ��NON ��PTB x�ESS h�ESB X�ESL D�ESO 0�ESC �ESD �ESF �ESE ܶESG ȶESH ��ESM ��ESN ��ESI ��ESA p�ESZ `�ESR L�ESU <�ESY (�ESV �SVF �DES �ENG �ENU �ENU ��USA ��GBR �CHN �CZE ܵGBR ̵GBR ĵNLD ��HKG ��NZL ��NZL ��CHN ��CHN ��PRI |�SVK l�ZAF `�KOR P�ZAF D�KOR 0�TTO �GBR  �GBR �USA �USA 6-0   OCP ACP Norwegian-Nynorsk   c c s   U T F - 8   U T F - 1 6 L E     U N I C O D E    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   ->* &   +   -   --  ++  ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        ������������|�t�h�\���������`�D�T�L�d�H�D�@�<�8�4�(�$��� ��������ȝ�� �������ĝ������������������������������������x�l�X�8����������x�T�4����ܿԿĿ������|�`�@���Ⱦ����\�8���Ľ��GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    1#QNAN  1#INF   1#IND   1#SNAN  CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           \�`�   RSDSk�+NL�qL�)�����:   C:\Program Files\MAXON\CINEMA 4D R13\plugins\Applink_Cinema4D\obj\Applink_Cinema4DR13_Win32_Release.pdb             �T�           d�p���    �       ����    @   T� �        ����    @   ��           ����                @���           �����    @�       ����    @   ��\�        ����    @   (�           8��                x�T�           d�l�    x�        ����    @   T�           ����l�    ��       ����    @   ��           ����l�    ��       ����    @   ��            ���           �(�D�    ��       ����    @   ���       ����    @   `�           p�x�    ��        ����    @   `�           ���           ������@�\�    �       ����    @   ��L�              P   �           �$�(�D�    L�       ����    @   ���              @   ���              @   `�            L��            ����           ������l�    ��       ����    @   ��            ����            ��    ��        ����    @   ��            ��8�           H�T��    ��       ����    @   8�            0���           ������l�    0�       ����    @   ��    P       P���           ��������@�\�    P�       ����    @   ��            ��,�           <�H��    ��       ����    @   ,�            ��x�           �����    ��       ����    @   x�             ���           �����     �       ����    @   ��             ��            �0����     �       ����    @   �            @�`�           p������    @�       ����    @   `�    X       ����           ��������@�\�    ��       ����    @   ��           ��,�    ��       ����    @   ����        ����    @   H�           X�,�                ��t�           �����,�    ��       ����    @   t�             ���           ����     �        ����    @   ��            <��           �(���    <�       ����    @   �             ���            x�l�           |�����    x�       ����    @   l�            ����           ����    ��        ����    @   ��            �� �           ����    ��       ����    @    �            ��L�           \�l����    ��       ����    @   L�           ����    �        ����    @   ��            ,���           ����    ,�        ����    @   ��            D��           (�4���    D�       ����    @   �            ��H�            ��x�           ����    ��        ����    @   x�            ����           ����    ��        ����    @   ��            ���           � �    ��        ����    @   �            ��P�           `�l���    ��       ����    @   P�            ���           ����    �        ����    @   ��            @���           �� �l�    @�       ����    @   ��            p�0�           @�P����    p�       ����    @   0�            D���           ����    D�        ����    @   ��            \�(�            d���           �����    d�       ����    @   ��            � (�           8�D��    �        ����    @   (�T ^  � \ �( �� �� ��  �  � @� `� �� �� Њ ��  � @� `� �� �� Ћ �� � 6� d� �� �� ό                         ��     ��   � �    @�    ����       ��     \�    ����       �            �	����    ����                  <�"�   L�   \�                            s            ����    ����                  "�   ��   ��                            ��              ��            �����    ����                   �"�   0�   @�                            ����    ����                  x�"�   ��   ��                            �����    ����                  ��"�   ��   ��                    �$    8�   H�d� �     �    ����    (   �-    ��    ����    (    -    c    ��   �� �    d�    ����       F            1����    ����                  ��"�   ��   ��                    �%     �   0�L� �    @�    ����    (   02     �    ����    (   �1            !6            6����    ����    ����    ����    "�   ��   ��                              x�            h�            �9            �8����    ����    ����    ����    "�   �   X�                              �            ��            �;            �;����    ����    ����    ����    "�   ��   ��                              ��            ��            �>����    ����                  �"�   �   ,�                            �D����    ����                  d�"�   t�   ��                            G����    ����                  ��"�   ��   ��                            �K����    ����                  �"�   $�   4�                            �M����    ����                  l�"�   |�   ��                            wR            wQ����    ����    ����    ����    "�   ��   (�                              ��            ��            �a����    ����                  P�"�   `�   p�                            �b����    ����                  ��"�   ��   ��                            �g            �g����    ����    ����    ����    "�    �   d�                              �             ������"�   ��                       ����.�"�   ��                       ����Q�    Y�"�   ��                       �����    ��"�   �                       ������"�   L�                           	    ��   ��d� �    p�    ����    (   �	    ����    ����    ����    Y    ����    ����    ����    p    ����    ����    ����    |    ����    ����    ����    �     ����    ����    ����    k"        7"����    ����    ����    �"    ����    ����    ����    �#    ����    ����    ����    �%    ����    ����    ����    %'    ����    ����    ����    \(    ����    ����    ����+,<,    ����    ����    ����    �.    ����    ����    ����    4    ����    ����    ����    _F    ����    ����    ����    �R        �R        �R    ����    ����    ����    �S    ����    ����    ����    �W    ����    ����    ����    �Z    ����    ����    ����    �^    ����    ����    ����    Qa����    `a����    ����    ����    c����    c����    ����    ����h!h    ����    ����    ����    �w    ����    ����    ����    d�    &�0�����    ����    ������@           �����    ����                  �"�   �   ,�                   ����    ����    ����    ,�    ��������    ����    ������    ����    ����    ��������    ʄ    ��   �� �    �     ����       b�    ����    ����    ��������    ����    ����    ����Ցّ    ����    ����    ����i�m�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    Z�    ����    ����    ����    ��    ����    ����    ����    3�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    
�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    !�    ����    ����    ����    �    ����    ����    ����'+'    ����    ����    ����{(�(    ����    ����    ����    �*    ����    ����    ����    K1    ����    ����    ����    �2    ����    ����    ����    ]7    ����    ����    ����    #9        _8����    ����    �����F�F    ����    ����    ����    �_H�          �  � ��          � T�                     �� �� �� �� �� ,� D� \� d� �� �� �� �� �� �� � *� >� P� `� l� x� �� �� �� �� �� �� �� � � � (� :� N� `� n� z� �� �� �� �� �� �� �� �� �� �  � .� @� L� \� n� �� �� �� �� �� �� �� � *� D� T� j� �� �� �� �� �� �� �� � *� :� P� `� p� �� �� �� �� ��     �     C CloseHandle EProcess32Next Module32First CProcess32First  � CreateToolhelp32Snapshot  KERNEL32.dll  ShellExecuteExA SHELL32.dll �InterlockedIncrement  �InterlockedDecrement  !Sleep �InitializeCriticalSection � DeleteCriticalSection � EnterCriticalSection  �LeaveCriticalSection  -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent ZRaiseException  �GetLastError  �HeapFree  �RtlUnwind � DeleteFileA �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �LCMapStringA  zWideCharToMultiByte MultiByteToWideChar �LCMapStringW  [GetCPInfo RGetACP  GetOEMCP  �IsValidCodePage �GetModuleHandleW   GetProcAddress  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �SetLastError  �GetModuleHandleA  �HeapCreate  �HeapDestroy WVirtualFree TVirtualAlloc  �HeapReAlloc �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA �WriteFile �GetConsoleCP  �GetConsoleMode  AFlushFileBuffers  hReadFile  �SetFilePointer  �GetModuleFileNameA  ExitProcess JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW �GetEnvironmentStringsW  TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �HeapSize  �GetLocaleInfoA  =GetStringTypeA  @GetStringTypeW  mGetUserDefaultLCID  � EnumSystemLocalesA  �IsValidLocale �InitializeCriticalSectionAndSpinCount �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW �SetStdHandle  �LoadLibraryA  �GetLocaleInfoW   CreateFileW x CreateFileA �SetEndOfFile  #GetProcessHeap      {qP    �          �� ��  � �� �   Applink_Cinema4DR13.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ̑��    .?AVApplinkDialog@@ ��    .?AVGeDialog@@  ̑̑��    .?AVbad_alloc@std@@ ��    .?AVexception@std@@ ��    .?AVfacet@locale@std@@  ��    .?AVcodecvt_base@std@@  ��    .?AUctype_base@std@@    ��    .?AVios_base@std@@  ��    .?AV?$_Iosb@H@std@@ ��    .?AV?$basic_istream@DU?$char_traits@D@std@@@std@@   ��    .?AV?$basic_ios@DU?$char_traits@D@std@@@std@@   ��    .?AV?$ctype@D@std@@ ��    .?AV?$basic_streambuf@DU?$char_traits@D@std@@@std@@     ��    .?AV?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    ��    .?AV?$codecvt@DDH@std@@ ��    .?AV?$basic_istringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    ��    .?AV?$basic_filebuf@DU?$char_traits@D@std@@@std@@   ��    .?AVlogic_error@std@@   ��    .?AVruntime_error@std@@ ��    .?AVlength_error@std@@  ��    .?AVfailure@ios_base@std@@  ��    .?AVbad_cast@std@@  ��    .?AV?$basic_ifstream@DU?$char_traits@D@std@@@std@@  ̑̑��    .?AVCommandData@@   ��    .?AVBaseData@@  ��    .?AVApplinkPreferences@@    ̑��    .?AVTriangulator@@  ��    .?AVCTriangulator@TRIANGULATOR@@    ̑̑̑̑��    .?AVGeModalDialog@@ ��    .?AVGeUserArea@@    ��    .?AVSubDialog@@ ��    .?AViCustomGui@@    ̑̑̑̑̑̑̑̑̑̑��    .?AVGeSortAndSearch@@   ��    .?AVNeighbor@@  ��    .?AVDisjointNgonMesh@@  ̑̑̑̑̑̑̑̑̑��    .?AVC4DThread@@ ̑̑̑̑̑̑��    .?AVGeToolNode2D@@  ��    .?AVGeToolDynArray@@    ��    .?AVGeToolDynArraySort@@    ��    .?AVGeToolList2D@@  ̑����̑��    .?AV_Locimp@locale@std@@    ̑   ̑��    .?AVout_of_range@std@@  ̑��8�8�<�@�H�H�P�X�`�h�p�x���    ̑
   Copyright (c) 1992-2004 by P.J. Plauger, licensed by Dinkumware, Ltd. ALL RIGHTS RESERVED.              ̑��    .?AVtype_info@@ N�@���D            u�  s�          ̑            fmod         D4F���F���F���F��������F�F���F�sqrt    H�J�   L�        ̑                                                                                                                                                                                                                                                                                                                                                abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     ��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����    C                                                                                              8�            8�            8�            8�            8�                                       H�ЧP�@@�   @����������                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 o&o&o&o&o&o&o&o&o&o&                                                                                                                                                                                                                                                                                         ̑��    .?AVbad_exception@std@@             `    `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����
                                                             p�   D�	   �
   ��   T�   $�    �   ԯ   ��   t�   <�   �   ܮ   ��   X�     �!   (�"   ��x   t�y   d�z   T��   P��   @���      x   
   ?         ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      ������������������������������*�>�N�n�s���������������1�6�V�j����������������&�:�Z�_�y�~�������������"�B�V�n����������������  ��� ���������ܴдĴ����������������������������x�l�d�\���T�L�D�8�0�$�������	         @.   ����������    .       �                                                                                                                                                                                                                                   �&         `�   d�   T�   X�   0�   (�!    �   L�   D�   4�   �   �   �   �    �   ,�   $�   �   �    �   ��   ��   ��   ��"   ��#   ��$   ��%   ��&   ��      �      ���������              �       �D        � 0     H�8�    �p     ����    PST                                                             PDT                                                             �	�	����        ����           ���5      @   �  �   ����             ������������   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l           �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                       �   0040E0t0�0�0�01H1z1d2�2;3�3�3�3�3�34434D4V4j4�4�4�4�4�6q7�7�7�788}8�8�8�8�8�8�899+9?9R9e9y9�9�9�9�9�9�9�9j:�:�:�:;M;_;�;�;�;<><k<�<�<=5=b=�=�=�=n>�>?!?2?H?R?�?�?      �   *0<0M0^0p0�0�0�0�0�0)1<1L1[1�1�1�1�1�12*2[2�4�4�45#5D5t5�5�56*6=6R6t6�6�67"7B7S7a7i7�7�78r8�8�8�8I9}9�9:<:g:�:�:�:�:;7;K;];f;};�;�;�;d<|<�<�<�<�<�<= =8=Q=i=�=�=�=�=�=>(>=>\>t>�>�>�>�>�>�>? ?$?(?,?0?4?8?<?@?D?H? 0  <  j2�2�2�2�2�2�233/3H3\3�3�3�3�3�3�3�3�344(4@4L4y4�4�4�4�4�45+5V5l5�5�5�5�5�5�566,6E6Z6r6�6�6�6�6�6�67,7C7b7w7�7�7�7�7�788-8?8Q8e8z8�8�8�8�8�8�8+9<9N9W9i9{9�9�9�9�9�9�9::.:@:U:i:�:�:�:�:�:�:�:;-;Z;t;�;�;�;�;�;�;<!<9<N<x<�<�<�<�<�<�<�<==$=<=H==�=�=�=�=	>">E>d>|>�>�>�>�>�>?%?@?W?v?�?�?�?�?�?   @  d  0#0B0W0r0�0�0�0�0�01'1;1P1e1y1�1�1�1�1�1�1
2272R2r2�2�2�2�2�2�2�23	3363P3o3�3�3�3�3�34.4\4s4�4�4�4�4�4�45%5<5[5p5�5�5�5�5�56'6<6W6n6�6�6�6�6�67 757J7^7s7�7�7�7�7�7�78818O8c8x8�8�8�8�8�8�8�8�899T9k9�9�9�9�9�9:>:S:i:}:�:�:�:�:�:;*;I;^;y;�;�;�;�;�;<*<E<\<{<�<�<�<�<�<=#=8=L=a=v=�=�=�=�=�=�=
>">O>a>s>|>�>�>�>�>�>�>�>??E?Z?r?�?�?�?�? P  d  0*0A0V0k0}0�0�0�0�0�011/1G1^1}1�1�1�1�1�12'2F2[2v2�2�2�2�2�2 33&383L3a3v3�3�3�3�3�34#454>4O4a4j4�4�4�4�4�4�4�45'5<5P5i55�5�5�5�5�5�56J6k6�6�677)7C7U7g7y7�7�7�7�7 88#8C8U8i8�8�8�8�8�8�899D9W9i9z9�9�9�9::%:.:?:Q:�:�:�:�:�:�:�:;.;I;^;g;y;�;�;�;�;</<A<J<[<m<�<�<�<�<�<==:=V=j==�=�=�=�=�=>>8>\>r>�>�>�>�>�>?$?6?>?R?k?�?�?�?�?�?�? `  H  0=0O0a0j0~0�0�0�0�01 1)1:1L1U1o1�1�1�1�1�1�1�12&2:2S2i2z2�2�2�2�2�2�23$3D3a3s3|3�3�3�3�3�3	44$454G4P4b4t485N5e5z5�5�5�5�5�5�566+6@6X6�6�677'797j7|7�7�7�7�7�7�78(8?8Q8e8z8�8�8�89T9f9�9�9�9�9�9r:�:�:�:�:�:�:�:;;.;B;Y;k;�;�;�;�;�;�;�;</<L<`<u<~<�<�<�<�<==L=`=o=�=�=�=�=�=�=>->>>P>Y>n>�>�>�>�>�>�>�>?%?M?�? p  �   80J00�0�0�0�0.1@1T1�1�1�1�1)2S2|2�2�23l3�3�344V4g4}4�4�4�4�45)5L5^5�5�5�5�56%6:6L6�6�6�6�6O7]7x7�7�7�7�7858C8P8�8�8�8�8�8$9E9i9�9�9�9�9�9::?:S:h:q:�:�:�:2;�;�;�;<�<�<�<==$=-=M=_=�=�=>+>�>�>�>�>�? �  t   �3�3�4n7�7�78+888z8�8�8�8�89G9m99�9�9�9�9�9�9�9
:!:;:P:l:�:�:�:�:�:;1;W;i;z;�;�;<�<�<�=�=5>J>�>�>?�?   �  x   	00d0u0�0�0�1�1�1,363[3�4�4�5�5�5�6�67�7�7�78�8�8�9L:�:@;S;m;�;�;�;�;<#<G<�<
=3=�=�=�=�=>5>�>�>??E?u?�?�? �  �   0!030n0�0�01T1�1�1�1'2A2S2�2�2�2(3t3�3�3494o4�4�4�4525U5�5�5;6y6�6�6
797�7�7�7�7u8�8�8<9\9v9�9�9�9�9�9�9::3:G:c:z:�:�:�:�:�:;;/;E;[;p;�;�;�;�;�;<$<=<�>�>�>?%?-?C?Z?v?�?�?�?�?�?   �  �   0k0�0�0	1e1�1�1�1�1�1�12262M2l2�2�2�2�2"3N3�3�34;4�5U6�6�6�6�6�7�7�8�89"919�9�9�9�9�9�9E:Y:n:�:�:�:�:�:;$;-;A;V;�;�;�;�;�;y<�<�<�<,=G=�=�=>L>h>�>�>?)?j?�?�?�?   �  �   $0@0^0�0�01�1�1�1�1L2g2|2�2�2�2�23"363K3`3�3�3�3�344.4x4�4�4�4�4V5k5�5�5>6�6�6�647j7�7�78?8�8p9�9�9�9�9�9�9�9::O:c:x:�:�:�:�:Z<�<�<�<�<==(=<=�=�=�=�=�=>1>F>Z>n>�>5?�?   �  �   �0�2�2�2�2�213�3�3�3�3 454J4�5�5�5616L6c6�6�6�67J7'8<8P8X8m8�8�8�8�899.9C9q9�9�9�9�9�9::!:t:�:�:�:�:�:;*;>;S;�;�;W<m<�=�=>>�>5?�?�?�?   �  x   i0q0|0�0�0�011S1�1�1�1�3$4�6�7A8�8_9�9�9�9b:�:�:�;�;�;<0<J<y<�<�<�<= =7=`=�=�=�=(>E>�>�>�>�>�>
?T?i?~?�?�?�?   �  �   00030H0�0�0�0�0�0�1�1�1�1�1�1�1�1T2i2}2�2�2D3q4�4�4�4�455.5B5W5y5�6�6�7�7�7�78!878L8�9�9�9�9I:T:�:�:�:�:�;�;�;�;�<�>�>�?�?   0   51�12@2�233L3�3�3N5Y5M669F9n;w;�;�;�?  (   �01�1&363�3�3^4�42566H6�687W;W?   D   �34R4q4�4�5�5�5G6�:�;�<=L=z=�=�=�=�=>>1>9>?>D>U>�>�>�>�? 0 P   �0�0o1�1�1�1�1�1	2I2g23-3f4x4V7k7�:�:==!=)=/=4=E=�=�=�=&>8>?)?;?f?�? @ <   ]2�3�3�56(647%9,989�9�9�9�9�9�9X:v:�:�;�;<�=�?�?   P 0   $6A6M6W6�6�6�6 77 727|7�7}9�:d;y;x<%>0> ` X   v1�1f2v2�56(=.=4=:=G=T=�=�=�=�=�=�=>>4>E>S>q>�>�>�>�>??4?L?`?p?�?�?�?�?�?�? p   040L0`0o00�0�0�011$1D1d1�1�1�1�1�12$2T2t2�2�2�2�23A3T3�3�3�3�3�3444Q4a4q4�4�4�4�45$5D5d5�5�5�5�5�56D6^6u6g7�7�7�7�7�7�7�8�8�8�89D9d9�9�9�9�9:$:D:a:t:�:�:�:�:;1;D;_;m;{;�;�;�;�;�; <!<D<d<�<�<�<�<�<�<�<=/===K=Z=l=�=�=�=�=>4>T>t>�>�>�> ??-?W?i?�?�?�?�?�?   �   040T0t0�0�0�0�0�0�0141N1b1q1�1�1�1�1�12,2=2K2b2w2�2�2�2�2�233&3t3�3�3�3�3444A4Q4d4�4�4�4�45$5D5d5�5�5�5�56$6D6d6�6�6�6�67$7D7d7�7�7�78$8D8d8�8�8�8�89$9D9d9�9�9�9�9:$:D:d:�:�:�:�:;$;D;a;t;�;�;�;�;<!<1<A<T<t<�<�<�<�<=$=I=j=�=�=�=�>�>??-?`?u?�?�? � �   040Q0d0�0�0�0�01D1t1�1�1�1�1�2�2�2343w3�3�4�4�4�4�4�4515Q5�5�5�56q6�6�6
7,7j7�7�7�7�7K8�8�8 909`9�9�9�9�9:.:G:v:�:�:�:;6;R;q;�;�;�;<%<P<o<�<�<�<=5=G=�=�=�=>$>K>]>�>�>�>??j?�?�?�?   � �   0�0�0;1�1�12=2h2�2�23I3c3�3�34K4v4�4�45.5T5�56�6�6%7d7�7�7�7=8�8�89a9�9�9�92:k:�:�:�:�:�:1;j;�;�;t<�<=`=�=�=@>�>�>S?�?   � �   0S0�01s1�132�2�2S3�34c4�4#5�5�56�6�6@7p7�7�7 808`8�8�8 9M9q9�9�9�9:N:�:�:
;[;�;�;><~<�<�<"=D=�=�=�=$>d>�>�>?5?N?t?�?   � �   E0J0U0k0�0�0141n1@2�233 3$3(3,3034383f34p4t4x4|4�4�4�4�4�465X5b5�5�5�5�56!6A6a6�6�6�67$7D7t7�7�7$8D8t8�8�8�8�9�9�9:1:Q:t:�:�:;4;Y;v;�;�;�;�;�;�;<$<B<`<q<�<�<�<�<�<�<==4=d=�=�=>$>T>�>�>�>$?d?|?�?�? � �   $0d0�0�0�0�1�12%2>2e2�23/3H3b374t4�45
55*5H5R5t5�5646T6v6�6�6�6�67�7�7U8�8�8949d9�9�9s:�:�:�:;1;q;�;�;�;�;<D<�<�<�<�<�<�<"=T=�=�>�>�>�>?2?E?e?�?�?�?�? � �   0,0j0�0�0�0+1?1Q1b1�1�1�1�12)272D2o2�2�2�2�2-3N3�3�3�3H4�4
5'5T5�5�5�566b6�6�67727K7]7y7�7�7�7�788,848G8_8t8�8�8�8�8�8�89$9;�;�;D<�<�<i=�=�=d>�>�>?�?�?   � �   x0�0D1]1�1�1�1�1�1�1(2I2f2�2�23-3@3L3�3�3�3�3�3"4>4m4{4�4�5�5;6E6�6�6�6717_7�7�7�7�78�8�8�89y9�9�9:y:�:�:�:�:;4;U;�;�;Q<�<�<?=T=t=�=�=�=�=>$>Q>t>�>�>�>�>?4?a?t?�?�?   �   0!0A0a0�0�0�0111Q1t1�1�12!2D2d2�2�2�2�23$3D3d3�3�3�3�3�3444�4�4�4L5w5�5�5Q6�6�67�7�7�7A8^8v8�89#9�9�9�9!:D:�:3;\;�;<,<T<�<�<$=�=�=�=K>�>�>A?g?�?�?    �   A0g0�0,1�1�1�1n2�2�23>3S3�3�34|4�4545Q5a5t5�5�5�56$6T6t6�6�6�6747Q7t7�7�78 8B8~8�8�8�899Q9q9�9�9�9�9�:�:�:�:�:�:;4;Q;d;�;�;�;�;<D<t<�<�<�<�<�<=4=W=�=�=�='>b>�>�>�>?$?Q?d?�?�?�?   �   0$0T0�0�0�0141T1�1�1�1�12$2D2d2�2�2�2�2�2�23$3D3d3�3�3�3�3$4D4d4�4�4�4�4�45545T5t5�5�5�5�5$6D6d6�6�6�6�6�67A7T7t7�7�7848T8t8�8�8�8�8949T9t9�9�94:c:�:�:4;a;�;�;�;<<D<d<�<�<�<�<�<=$=D=y=�=�=>%>H>t>�>�>�>?&?6?d?�?�?�?�?�? 0 �   040T0t0�0�0�0�0121T1z1�1�1�1�12222B2d2~2�2�2�2�23/3T3l3�3�3�3�3�3$4<4e4�4�4�4�4�45K5^5�5�5�5�546T6t6�6�6�67$7D7d7�7�7�7�7�7$8D8d8�8�8�8�89$9D9d9�9�9�9�9�9�9$:A:T:q:�:�:�:�:�:�:;�;<B<u<�<�<%=u=�=�=>E>�>�>
?Q?�?�?   @ �   0U0�0�0�0E1�1�12U2�2�2�253r3�3�3%4u4�4�455x5�5�5�5�56U6�6�67U7�7�728�8�8�8�890959]9�9�9�9�95:Y:�:�:;9;b;�;�;�;<X<�<�<�<)=x=�=U>r>�>�>�>�>?$?D?a?q?�?�?�?�?�?�?   P �   040T0t0�0�0�0�0111T1�1�1�1�12$2D2d2�2�2�2�23$3D3a33�3�3�3�3$4O4q4�4�4�4�4515D5d5�5�5�5�5�5$6D6d6�6�6�6747a7�7�7�78d8�8�8949T9t9�9�9�9�9$:4:d:�:�:�:;$;T;t;�;�;�;<O<q<�<�<�<'=Q=q=�=�=�=�=>1>Q>q>�>�>�>�>?1?Q?q?�?�?�?   ` �   00D0d0�0�0�0�01!1A1T1�1�1�1�12!2D2d2�2�2�2�2313T3t3�3�3D4�4�45$5D5d5�5�5�56$6Q6t6�6�6�6$7Q7t7�78!8A8d8�8�8�89!9A9a9�9�9�9:4:Q:t:�:�:�:;1;T;q;�;�;�;�;<d<�<�<=$=Q=t=�=�=�=!>D>q>�>�>�>�>A?d?�?�?�?   p �   040d0�0�0+1T1�1�1�1�12A2d2r2w2�2�2�23j3�3�3�3$4D4�4�445�5�5�5
6-6a6�6�6�67/7t7�7�7�78I8�89$9Q9t9�9�9::5:T:�:�:�:�:;4;d;�;�;�;�;1<T<�<�<�<�<=4=q=�=�=�=A>d>�>�>�>?.?J?f?�?�?�? � |   0A0a0�0�0�0�0�0&1H1^1v1�1�1�122W2u2�2�2�2�2303L344R4e4�4�4�45+7�9�9D:W:�:�:�:;/;�<�<�<�<[=`=�=�=E>�>?U?�?�? � �   40d0�0$1X1�1�1�1�1�1$2V2�2�2�2�2�2&3;3Y3u3�3�3�3�3484m4{4�4�4�455*5G5t5�5�7k8�8�8�8+9f9�9�9�9�9�9�9::&:9:K:]:o:x:�:�:�:�:�:;%;8;d;r;;�;�;�;�;�;�;<$<6<R<h<�<�<�<�<�<�<="=3=F=t=�=�=�=�=�=�=�=�=>4>F>b>x>�>�>�>�>�> ??2?D?V?_?}?�?�?�? � �   00070I0[0m00�0�0�0�0�01$161H1Q1o1�1�1�1�1�1�12.2D2b2o2�2�2�2�2�23D3a3�3�3�344 4;4W4p4�4�4�4�4565X5u5�5�566$6}6�6�6�6�6�6727O7�7�748I8k8�89919A9T9�9�9�9�9�9:4:Q:d:�:�:;<< <'<.<5<<<C<J<x<�<�<}=�=z?�?�?   � �   0�0�0�0�0�0�0�0�0�0�0�0�0�0�01	11�2�2�2�2�2�2�23.3b3u3�3�3�3�3�3�3�3�3�3474�45E5\5q5z5�5�56&646z6�6�6747Q77�7�7E8Q8[8a8f8�8�8�8�8919D9a9t9�9�9�9::#:(:T:k:�:�:�:!;A;a;�;�;   �    6   � p   a0�0�0�0%1e1�1�152r2�2�23R3�3�34E4�4�4�45B5u5�5�5E6�6�67U7�7�7E8�8�859u9�9�;�;^>�>�>�>�>�>�?�?�?�?   � �   �0�0�0�0~1�1�1�1�123*3C3Q3�3�3�3�3�4�4�45!545d5�5�5�5�5646d6�6�6�67$7D7a7t7�7�78(878t8�8�8�8919T9t9�9�9�9:1:�:�:�:4;Q;d;x=�=�=�=�>�> � t   (0a0t0�0�0�0!111A1Q1s1�1�1�1242W2e2t2�2�2�23!343d3�3x4�4
55{5C6V6f677&7�7�7�7Q8t8�89D9�9�9z=>>L?�?�?   �   0060U0f0�0�0-1�2�233 3&303?3^3{3	44%41494?4N4W4�4�4�4�45!5R5y5�5�5�5�5�566\6i6s6x6�6�6r7{799!9A9K9h9y9�9�9�9::-:N:�:�:�:
;;&;9;@;K;Q;\;a;�;�<�<�<�<�<�>�?�?  �   0!0'0+01050;0?0E0I0N0T0X0^0b0h0l0r0v0�0�0�011'1,10141]1�1�1�1�1�1�1�1�1�1�12222 2�2�2�2�2�2�2�2�23=3D3H3L3P3T3X3\3`3�3�3�3�3�3P4d4�45#5;5X5e5�5S7e778A8N8i8p8�8�8�899g9m9~9�9�:�:�: =@=z=�=�=>>~>�>�>??�?�?�?   p   {0�1�1�1�1=2w2�2�335�6�7q8{89�9[:`:j:�:�:�:�:
;;+;[;w;�;�;<�<�<�<g=�=�=�=�=�=^>p>�>�>�>?.?�?�?�?�?   0 �   0000=0c0�0�0�0�0�0�0�0�0�0�0�0�0�0 1f1q1�1�1�1�1�1�1�12$2(2,2024282<2@2�2�2�2�2�2�2�2u3�3�3�3�314;4H4�4�455535E5R5^5h5p5{5�5�5r6"7E7�7�8 9(9�9�9: :�:�:;#;�;�;�;�<T>?.?8?B?m?u?�?�?�?�?�? @ �   00(0a0j0v0�0�0�0w1�1�1i2v2�2�2�2�283�3'4r4�45U5�5�5	6E6l6u6~6�6�6�6�6�6f78_8�8�8�8�8�8T9m9~9�9 :�:�;Q<4>d>�>�>?S?�?�?   P �   30;0e1	22M2W2c2l2�2Z3R4g45A7a7f7�8�8�8a:r:�:�:�:�:�:�:;#;-;F;P;c;�;�;�;<v<�<�<G=f=�=�=�=>'>/>7>N>g>�>�>�>�>�>�>�>�>?#?)?4?@?U?\?p?w?�?�?�?�?�?�?�?�?   ` �   
000(070=0F0R0`0f0r0x0�0�0�0�0�0�0�0�0	1/1o1u1�1�1�1�1�1y2�2�2�2�223B3H3T3Z3j3p3�3�3�3�3�3�3�3�3�3�3�3�3�3�34	444#4(4.42484=4C4H4W4m4x4}4�4�4�4�4�4�4�4�4�4�45P5l5�5�56666 6&6-646;6B6I6P6W6_6g6o6{6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�7�84;�;�; p �   +1�1�3�3�3444#4�5�5�5�5�5�5�5�5666'6/696?6E6R6Y6c6�6�6�6�6�6�6�6�677>7�7�788I:W:]:w:|:�:�:�:�:�:�:�:�:�:�:�:;;$;);1;7;A;H;\;c;i;w;~;�;�;�;�;�;�;�;�;F<�?�?   � @   !0G0�0�0�2�2�2�2�22344,4D4�4�4�4�4�5�6�78�9*;B>i>v>   � �   t0h1�1�1�1�1M2S2m2|2�2�2�2�2�2�2�2�2
33-373]3�3�3�3�3�3�4�4/5C5d5j5�5�5�5;6E6m6�6�6�6	7[7a7�7�7�799k9�9":�:�:�;<h<�=�>�?�?�? � P   '0F0�01F1�1�12J2T2�2=34�46�6�6�6�67?7>8�8�9T:�:�:�:�:;?;|<�<=A=   � ,   #4o>v>�>�>�>�>?%?,?5?u?z?�?�?�?�?   �   0)0M0w0�0�1�1�122=2X2^2g2n2�2�2�2
333*343;3F3O3e3p3�3�3�3�3�344:4?4J4O4m4�4555U5_5�5�5�5�5�5�7�7�7�7�7�7)8/8E8P8g8s8�8�8�89 9R9k9z99�9�9�9V:\:u:{:K;n;{;�;�;�;�;�;�;<<<�<�<�<�<==&=2=W=`=i=v=�=�=�=�=�=�=�=�=�=>>>T>X>\>`>d>h>l>p>t>x>|>�>�>�>�>�>?z?�? � D   {0�0�0�041q1�1�2�2�2�2�2�2�304�4L5�5�5�5�5�5h6�6�=�>�>E?�?�? � �   0M0�1�1�1�2�2�2�3�4�4�4�4�4�4�45>5w5�5c6r6�7�7�7�7�7�7�7�7(8�869�9�9:W:]:i:�:�:);�;�;�;�;<8<l<r<~<�<Z=_=d=i=y=�=�=�=>G>L>S>X>_>d>�>�>�> � P   #55�5�5�5�577"7E7�7�7�7�7�788S8U:�:�:�<�<�<=I=Y=k==�=,>�>�>�>?     (   �0
1�1�122e2�2�2�23^3q3�3�3�8  p   :::#:':+:/:3:7:;:?:C:G:K:O:S:W:[:_:c:g:k:o:s:w:{::�:�:�:�:�:�:�<�<�<=t=�=�=�=�=
>7>?>^>n>�>�>�>�>�?   T   �12�2�4�6�67;7�7�78-8A8G8�819=9�9�9�9�9:':N:[:`:n:�:;�<M=W=>>�>�>v?�? 0 �   0[0�0�0�1�1�1�12J23E3`3n3v3�3�3�3�3�3�3�3�3�34�4%5]5p5�5�5�5�56,6�6�6�6�6E7P7~7�7�7�7�7I8V8~8�8�8�8�9�9�9�9::":1:7:F:L:Z:c:r:w:�:�:�:�:	;H;O;U;�;�;�;�;�;�;�;�;�<�<2=�?   @ D   /1J1`1v1~1�1�2b3�3�3F4W6i6{6�6�6�6�6�7d8�8�89969�<q=�>*?O? P H   21.32363:3>3B3F3J3l3`4�5�6�9U:�:�:�:;;&;f;�;i>�>�>�>	??+?P?g? ` D   0E1A2344�4�5I6O6�6�67�7�7a8W9_9:�:�;�;5<;<K<�<=2=�=   p 4   �0�0�3�3�3�344	444444*455-5Y5�5�5�? � �   �1�1�1�1�1�1�1�13&3<4C4�4�4!5N5�5q6\7x7�9�9�9�9�9:2:R::�:�:�:;2;R;r;�;�;�;<%<H<v<�<�<�<�<�<===)=5=B=J=T=f=p=�=�=�=�=�=   � �  `1d1h1l1p1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8�8�8$;(;,;0;4;8;<;@;D;H;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<0=4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=(>,>0>4>8>�>�>�?�?�?�?�?   � h   H0L0�0�0�0�0�0�0�0�0�0�0�0�1�1�1�1�1�1�1�1�1�1�1�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�;�; <$<(<,<   � �   : :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�< � l  �2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4�6�6L7P7`7d7h7p7�7�7�7�7�7�7�7�7�7�7�788$84888L8P8`8d8l8�8�8�8�8�8�8�8�8�8�8�89999 9(9@9D9\9l9p9x9�9�9�9�9�9�9�9�9�9�9�9 :::::$:<:@:X:\:t:�:�:�:�:�:�:�:�:�:�:�:�:�: ;; ;0;4;D;H;L;T;l;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<$<(<8<<<@<H<`<p<t<�<�<�<�<�<�<�<�<�<�<�<�<=== =$=(=0=H=X=\=l=p=t=x=�=�=�=�=�=�=�=�=�=�=�=�= >>>>(>,>D>T>X>l>p>�>�>�>�>�>�>�>�>�>�>�>�>???? ?(?@?P?T?d?h?x?|?�?�?�?�?�?�?�?�?�?�?�?   � �  000040D0H0X0\0`0d0l0�0�0�0�0�0�0�0�0�0�0 111$1(1,141L1\1`1p1t1�1�1�1�1�1�1�1�1�1�1 2222 282H2L2\2`2d2l2�2�2�2�2�2�2�2�2�2�2�2�2 33(3,3<3@3D3H3P3h3x3|3�3�3�3�3�3�3�3�3�3�3�3�34 4$44484<4D4\4�4�4�4 555$585H5l5x5�5�5�5�5�566,6P6\6d6�6�6�6�6�6 777,747<7@7D7L7`7h7|7�7�7�7�7�7�7�7�7�7�788$8(8,848H8P8d8t8�8�8�8�8�8 99<9D9h9|9�9�9�9�9�9::<:H:P:p:�:�:�:�:�:�: ; ;D;P;X;x;�;�;�;�;�;<<8<L<\<�<�<�<�<�<�<�<==H=P=t=�=�=�=�=�=�=�=�=>$>0>P>\>|>�>�>�>�>�>�>�>�>?0?P?\?x?�?�?�?�? � �   0080X0x0�0�0�0�0�0101P1\1x1�1�1�1�1�1�1�1222<2H2P2�2�2�2�2�2�2�2�2�2�2�2�2 33 3<3@3\3`3�3�3�3�3 4 4@4`4�4�4�4�4�4 55 5@5`5�5�5�5�5�5�56 � (   00 080<0@0\0x0�0�0�0�01L1�1�1�102P2�2�2 3 3@3d3�3�3�3�3�3�34 4<4h4l4p4t4x4�4�4�4�4�4�4�4�4�4�4 5555,5D5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5646<6@6d6l6p6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6@7D7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88<�=�=�=�=�=�=>>>>> >$>�?�?�?�?�?�?�?�?�?�?   p  �0�0 1(1�3�3�3�34444$4,444<4D4L4T4\4d4l4t4|4�4�4�4�4>5B5F5J5N5R5V5Z5^5b5f5j5n5r5v5z5~5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�566
666666"6&6*6.62666:6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$707l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89999$9,949<9D9L9�9�90:4:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            