MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       l���(���(���(��k�*���!�h�7���!�~����'��-���(���H���!�y�q���!�o�)���!�l�)���Rich(���                        PE  L ���N        � !	  Z  �      �     p                         `                              0� S   d� <                             �5  �q                            (� @            p \                          .text   �Y     Z                   `.rdata  �[   p  \   ^             @  @.data   ;   �     �             @  �.reloc  LA     B   �             @  B                                                                                                                                                                                                                                                                                                                                                                                        U��t�V��H�QV�ҡt��H�U�AVR�Ѓ���^]� U��t�V��H�QV�ҡt��U�H�E�IRj�PV�у���^]� ����������U��t��P�E���   ��VWP�EP�E�P�ҋu���t��H�QV�ҡt��H�QVW�ҡt��H�A�U�R�Ѓ�_��^��]� ������������V���X` �N��q�[ �N$�B9 ��^���������������V��N$��q�: �N��[ ��^�?` ���������������U���T  ��3ŉE�Wj j�8 ����u_�M�3���� ��]�V������PWǅ����(  �^8 ����   ������Qj�N8 �����   ������RPǅ����$  �"8 ���}   ������P������h  Q��� ������h  R�`� ���������P�I �@��u�+�$    ��/t��t������H��\uꍴ����V�5� hrV��� ����u.������PW�7 ���8���W� p^3�_�M�3���� ��]ËM�^3͸   _�� ��]���������j j j�Ń �����U���\V��E�P�M�Q���E�   �E�    �k �}� �  W�M��g7 �t��B�P�M�Q�҃��E�Pj�M܍~Q���n���P�M��7 �U�R�M��	; �M��8 �t��H�A�U�R�Ћt��Q�J�E�P�у�h�r�M��7 �U�R�M���: �M���7 �E�j P�?G �����M  �t��Q�J�E�SP�ыt��B�Pj j��M�h�rQ�ҍE�P�-� �t��Q�J�E�P�у�j ���` �t��B�P�M�Q�ҡt��H�Aj j��U�h�rR�ЍM�jQ�x� �t����B�P�M�Q���҃� j ����   hpr�M�������E�P�� �t��Q�J�E�P���� hrh�   h��h�   ���� ����t	���M�  �3�WS����  h�  ����_ [�M��6 _^��]� j �U�R���E�   �E�    般 [�M��_6 _^��]� �������U���SVW��j�~W�E�3�P�E�   �]�芭 jW�M�Q���E�   �]��r� jW�U�R���E�   �]��j jW�E�P���E�   �]��Bj jW�M�Q���E�   �]��*j jW�U�R���E�   �]��j jW�E�P���E�   �]���i jW�M�Q���E�   �]���i j
W�U�R���E�
   �]��*j j	�E�	   �]�W�E�P���i jW�M�Q���E�   �]��i jW�U�R���E�   �]��i jW�E�P���E�   �]��j� jW�M�Q���E�   �]��Ri _^[��]������������U���   V���?� ��u^��]�SWh s�M���3 �E�P�M�Q�~$�H ��P�U�R��7 ��P���7 �M��4 �M��4 �M��w4 3ۉ^@��I SW�E���C ������  �E�P���5 P�M���3 jj�M�Q�M�htaoc��I ���M��E��!4 �t��B�P�M�Q�҃�8]�t�E�P�I ��_[3�^��]�Sh�r�M�������t��Q�R8�E�P�~j���ҡt��H�A�U�R�Ѓ�h�r�M���2 h�r�M���2 �M�Q�U�R��l���j	P��G ��P�M�Q��6 ��P�U�R��6 ���M��b3 ��l����W3 �M��O3 �M��G3 �E�jP�B ���M̅�t0Q�M���3 �t��RP�B8j���Ћt��Q�J�E�P���ZSh�r�����P�� �t��B�P�M�Q�҃�Sh�r�M�������t��P�R8�E�Pj���ҡt��H�A�U�R�Ћt��Q�B4��Sj���Ћt��Q�B0jj���Ћt��Q�B0jj���Ћt��Q�B0Sj���Ћt��Q�B0Sj���Ћt��Q�B0jj���Ћt��Q�B4Sj
���Ћt��Q�B0jj	���Ћt��Q�B0jj���Ћt��Q�B0Sj����Sh�r�M�������t��Q�E�Pj�ϋR8�ҡt��H�A�U�R�Ћt��Q�B0��Sj���ЋM�W��M �M��VG �M��~1 �M�Q�N$�22 P�M���0 �M�jj�U�Rhtaoc�G ���M��E��F1 �t��H�A�U�R�Ѓ�8]�t�M�Q�F ��_[3�^��]ËM�j�~W�I �M���F �t��E�   �]�B�P�M�Q�҃�SS�E�Pj�M�Q������P�U�R����` �t��H�A�U�R�Ћt��Q�J�E�P�ыt��E�   �]�B�P�M�Q�҃�SS�E�Pj�M�Q������P�U�R���` �t��H�A�U�R�Ћt��Q�J�E�P�у��E�   �]�h����t��B���   h  �Sjh���h  �Sj����P�E�P���:[ �t�S�E�   �]�Q���   Sj����P�M�Q���� �t�S�E�   �]�B���   Sj����P�E�P����� �t�S�E�   �]�Q���   Sj����P�M�Q��蓥 �t�S�E�   �]�B���   Sj����P�E�P���f� �t��E�   �]�S�Q���   Sj����P�M�Q���9� �t�h���h  �Sjh���h  ��E�
   �]�B���   Sj
����P�E�P���Z �t�S�E�	   �]�Q���   Sj	����P�M�Q���ɤ �t�S�E�   �]�B���   Sj����P�E�P��蜤 �t�S�E�   �]�Q���   Sj����P�M�Q���o� �t��E�   �]�B�M̋PQ�҃�SS�E�Pj�M�Q���]���P�U�R���1^ �t��H�A�U�R�Ћt��Q�J�E�P�ыt���S�E�   �]�B���   Sj����P�E�P���ޣ h�  ���W �M�Q�9C ��_[�   ^��]�����������U���0V��~@ t~W��B �E��E�P�N$�,. P�M���, jj�M�Q�M�htaoc�C �MЋ��D- �t��B�P�M�Q�҃���_t��������M���V�gI �M���B �E�P�B ��^��]���������������U���   SV��3�W�]��F@   �����E����   ����   ����  �t��H�A�U�R�Ћt��Q�JSj��E�hprP�эU�R�/� �t��H�A�U�R���I� hrh�   h��h�   ���.� ��,;�t�����  ��VW���D�  _^�C[��]� ��3�VW���*�  _^�   [��]� �MQ�U�R���E�   �]��^ 9]�1  h�  ���>U _^�   [��]� �� hrh�   h��j$��蓸 ��;�t�@   ��X�X�X�X�3���VW���gO  �t��H�A�U�R�Ѓ��M�Qj�U�R�������t��H�A�U�R�Ћt��Q���   ��Sj���Ѕ�t2Sh�r�M��&����t��Q�Rx�E�P�M��E�   ���E��u�]�E�t�t��H�A�U�R�Ѓ�8]�  ���������   �t��Q�Bdj�M��Ћt��Q�����   hrFh�   V�Ћt��Q��j���BhVW�M���j<��X���SQ�� ����X���RǅX���<   ��\�����`���ǅd���<s��h�����p���ǅt���   ��x����Tq��uVSh$s�M������E�P�� �t��Q�J�E�P���(Shs�M�������U�R�� �t��H�A�U�R�Ѓ��t��Q�J�E�P�у�_^�   [��]� �����������VW��3�9>t	V�p� ���>�~�~�~�~_^�������������U��V��N$��q�\) �N�4K ���O �Et	V�a� ����^]� �������U�������M�P�P�P�P �P(�P0�P8�P@�PH�PP�XX���Q�P�Q�P�Q�P�Q�P�I�H�M��P�Q�P�Q�P �Q�P$�Q�P(�I�H,�M��P0�Q�P4�Q�P8�Q�P<�Q�P@�I�HD�M��PH�Q�PL�Q�PP�Q�PT�Q�PX�I�H\]� �����������U��M�U�A�
�E��B�I0���B�IH����A �
�A�A8�J���AP�J���X�A(�
�A�A@�J���AX�J���X�A�J�B �I0���B(�IH���X�A8�J �A �J���AP�J(���X �A@�J �A(�J���AX�J(���X(�A�J0�A0�J8���AH�J@���X0�A8�J8�A �J0���AP�J@���X8�A@�J8�A(�J0���AX�J@���X@�A�JH�BP�I0���BX�IH���XH�BP�I8�BH�I ���AP�JX���XP�A@�JP�BH�I(���AX�JX���XX]���U��t��UV��H�AVR�Ѓ���^]� ��������������U��t��H�U�I(��VWR�E�P�ыt��u���B�HV�ыt��B�HVW�ыt��B�P�M�Q�҃�_��^��]���U��t��E�H�U �E��VWR�UP�ERP�A$���U��$R�Ћt��Q�u���BV�Ћt��Q�BVW�Ћt��Q�J�E�P�у�,_��^��]��������������U���$�ESVW3ۍM�Q�M��]܉]�E�]��]�� �}S�U�R�E�P���d	 �M����� ;�th�t����   �JX�E�P�ы���;�tJ�t����   �PT���ҋt��Q|�M�RQPV�ҋ�t����   ��U�R�Ѓ�_��^[��]� �t����   �
�E�P�у�_^3�[��]� ������������U���$�EVW3��M�Q�M��}܉}�E�}��}���  �MW�U�R�E�P� �M����� ;�tZ�t����   �JH�E�P�ыt��u���B�HV�ыt��B�HVW�ыt����   ��M�Q�҃�_��^��]� �t��H�u�QV�ҡt��H�QWj�h�rV�ҡt����   ��U�R�Ѓ�_��^��]� ��������U���$�EVW3��M�Q�M��}܉}�E�}��}���� �MW�U�R�E�P� �M������ ;�t8�t����   �J8�E�P�ыt������   ��M�Q�҃�_��^��]� �t����   ��U�R�Ѓ�_3�^��]� �U���$�ESV3��u��M�Q�M��u܉u�E�u��u��5� �MV�U�R�E�P�� ��t �t����   �J�E�P�у���t��2ۍM��� ^��[t7�t����   �P<�M�Q���]�t����   ��U�R���E����]� �t����   �
�E�P���E����]� ���������U���$�EVW3��M�Q�M��}܉}�E�}��}��h� �MW�U�R�E�P�' �M����]� ;�t[�t����   �J@�E�P�ыu��H��P�N�H�V�P�@�N�t��V���   �
�F�E�P�у�_��^��]� ��t��u����   �V��^�M�Q�҃�_��^��]� U���$�EVW3��M�Q�M��}܉}�E�}��}��� �MW�U�R�E�P�W �M����� ;�tD�t����   �JL�E�P�ыu��P���V! �t����   ��M�Q�҃�_��^��]� �uW���  �t����   ��U�R�Ѓ�_��^��]� ����������U��Q�t��P�BdVWj�M�Ћt��Q�����   hPsFh�  V�Ћt���j�E��QVP�Bh�M��N3���~S�]�I �M��R���+ G;�|�[�E�P袩 �t��Q�J�EP�у�_^��]� �����U����t��H�AV�U�WR�Ћt��Q�Jj j��E�h�sP�ыt��B�Pd��j�M��ҋ�t��H���   hPsFh�  V�ҋt���j�E��QVP�Bh�M���N3���~S�]���M��R����* G;�|�[�E�P�Ҩ �t��Q�J�E�P�у�_^��]� �����U��Q�ESVW���   3�3�3�3ۃ��M�|#�@|�O���A�	�d$ p����u�E�M�;�}�@|��_�^�[��]� �����U��t��H�Q��   V�uV�ҡt��H�Qj j�hLtV�ҋE����
�  �$��. j hHt�M������E�P���nc  �t��Q�J�E�P����  j hDt��`����������`���R���7c  ��`����  j h<t�M������M�Q���c  �t��B�P�M�Q���p  j h8t�M������E�P����b  �t��Q�J�E�P���?  j h4t�M��[����U�R���b  �U��  j h,t�M��9����M�Q���b  �t��B�P�M�Q����   j h(t�M������E�P���]b  �t��Q�J�E�P���   j h t�M�������U�R���,b  �U��   j ht�M������M�Q���
b  �t��B�P�M�Q���kj ht��p���������p���P����a  �t��Q�J��p���P���4j ht��P����M�����P���R���a  ��P����t��H�AR�Ѓ��t��Q�J�E�P�ыt��B�Pj j��M�htQ�ҡt��P�B<�����Ћt��Q�RLj�j��M�QP���ҡt��H�A�U�R�Ѓ���^��]� �I , 9, d, �, �, �, - J- l- �- �- ����S�   V3�W���7�G�w�w�w�w�G(�w�w�w,�w$�w �G@�w0�w4�wD�w<�w8�GX�wH�wL�w\�wT�wP�Gp�w`�wd�wt�wl�wh���   �wx�w|���   ���   ���   �_���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   97t	W舤 ���7�w�w�w�w93t	S�m� ���G0�3�s�s�s�s90t	P�O� ���GH�w0�w4�wD�w<�w890t	P�0� ���G`�wH�wL�w\�wT�wP90t	P�� ���Gx�w`�wd�wt�wl�wh90t	P�� �����   �wx�w|���   ���   ���   90t	P�ǣ �����   ���   ���   ���   ���   ���   90t	P薣 �����   ���   ���   ���   ���   ���   ��_^[����������SVW����� ���   3�93t	S�D� ���3�s�s�s�s9��   ���   t	S�� ���3�s�s�s�s9wx�_xt	S� � ���3�s�s�s�s9w`�_`t	S�� ���3�s�s�s�s9wH�_Ht	S�¢ ���3�s�s�s�s9w0�_0t	S裢 ���3�s�s�s�s9w�_t	S脢 ���3�s�s�s�s97t	W�i� ���7�w�w�w�w_^[�����U���  �t�SVW���H�A�U�R�}��Ћt��Q�Jj j��E�hltP�ыt��B�P�M�Q�ҡt��H�Aj j��U�h`tR�ЋU��(�M�QR�E�P����P�M�Q�U�R�d  ��P�E�P�d  �t��Q�J�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ы]��S�t��B�H����V�ыt��B�P�M�VQ�҃��������u�~ �E�    ��  3��t��H�A�U�R�Ћt��Q�Jj j��E�h�sP�ыt��B�P�M�Q�ҡt��H�Aj j��U�h\tR�Ћt��Q�J�E�P�ыt��B�Pj j��M�h\tQ�ҡt��H�A��8���R�Ћt��Q�J��@j j���8���hXtP�ыF�t��D8��j0j jǋB�P$j ���������$Q�ҋءt��H������AR�Ћt��Q�J�����PS�ыt��B�P������Q�ҋF�D8��,j0j ǡt��H�A$jj ���������$R�Ћt��Q�J�؍�(���P�ыt��B�P��(���QS�ҡt��H�A������R�ЋF�t��8�Q�J$��,j0j j�j ��������$P�ыt��؋B�P��H���Q�ҡt��H�A��H���RS�Ћt��Q�J�����P�ыt��B�P�M�Q�ҡt��H�I�U�R��8���P�ыt��B�P<��8�M��ҋt��Q�RLj�j���H���QP�M��ҡt��H�A�U�R�Ћt��Q�R�E�P�M�Q�ҡt��P�B<���M��Ћt��Q�RLj�j��M�QP�M��ҡt��H�A��h���R�Ћt��Q�R��h���P�M�Q�ҡt��P�B<����h����Ћt��Q�RLj�j���(���QP��h����ҡt��H�A�U�R�Ћt��Q�R�E�P��h���Q�ҡt��P�B<���M��Ћt��Q�RLj�j��M�QP�M��ҡt��H�A��x���R�Ћt��Q�R��x���P�M�Q�ҡt��P�B<����x����Ћt��Q�RLj�j������QP��x����ҡt��H�A��X���R�Ћt��Q�R��X���P��x���Q�ҡt��P�B<����X����Ћt��Q�RLj�j��M�QP��X����ҡt��H�I�U�R��X���P�ыt��B�P��X���Q�ҡt��H�A��x���R�Ћt��Q�J�E�P�ыt��B�P��h���Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P��H���Q�ҡt��H�A��(���R�Ћt��Q�J�����P�ыt��B�P��8���Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҋE�t��Q��<P�B����S�Ћt��Q�J�E�SP�ыM܃������E�@��;F�E��j����}܋]�t��B�P�M�Q�ҡt��H�Aj j��U�hltR�Ћt��Q�J�E�P�ыt��B�Pj j��M�hPtQ�ҡt��H�U�I(R�����P�ыt����B�P�M�Q�ҡt��H�A�U�RV�Ћt��Q�J�����P�ыt��B�P�M���@Q�ҡt��H�I�U�R�E�P�ыt��B�P<���M��ҋt��Q�RLj�j��M�QP�M��ҡt��H�A�U�R�Ћt��Q�R�E�P�M�Q�ҡt��P�B<���M��Ћt��Q�RLj�j��M�QP�M��ҡt��H�I�U�R�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt���S����Q�BV�Ћt��Q�J�E�VP�у����m���S�������t��B�P�M�Q�҃�_^[��]� �������U���  �t�SVW���H�A�U�R�}��Ћt��Q�Jj j��E�h�tP�ыt��B�P�M�Q�ҡt��H�Aj j��U�h`tR�Ћu�F,��(�M�QP�U�R����P�E�P�M�Q��[  ��P�U�R�[  �t��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�ЋM���t��BQ�H����S�ыt��B�P�M�SQ�҃����'���3�9]�]��  �t��H�A��(���R�Ћt��Q�Jj j���(���h�sP�ыt��B�P������Q�ҡt��H�Aj j�������h\tR�Ћt��Q�J������P�ыt��B�Pj j�������h\tQ�ҡt��H�A��h���R�Ћt��Q�J��@j j���h���h�tP�ыF�t���j0�<[�j �j��D8ǋB�P$j ���������$Q�҉E��t��H�A������R�Ћt��Q�M��R������PQ�ҡt��H�A������R����F�d8�t��Q�J$��,j0j �jj ���������$P�ыt��E��B�P������Q�ҡt��H�E��I������RP�ыt��B�P������Q�ҋF�8��,j0j ǡt��H�A$jj ���������$R�Ћt��Q�J�E���H���P�ыt��B�U��@��H���QR�Ћt��Q�J������P�ыt��B�P��8���Q�ҡt��H�I��8���R��h���P�ыt��B�P<��8��8����ҋt��Q�RLj�j���H���QP��8����ҡt��H�A��X���R�Ћt��Q�R��X���P��8���Q�ҡt��P�B<����X����Ћt��Q�RLj�j�������QP��X����ҡt��H�A��x���R�Ћt��Q�R��x���P��X���Q�ҡt��P�B<����x����Ћt��Q�RLj�j�������QP��x����ҡt��H�A������R�Ћt��Q�R������P��x���Q�ҡt��P�B<���������Ћt��Q�RLj�j�������QP�������ҡt��H�A������R�Ћt��Q�R������P������Q�ҡt��P�B<���������Ћt��Qj�j�������QP�RL�������ҡt��H�A������R�Ћt��Q�R������P������Q�ҡt��P�B<���������Ћt��Q�RLj�j���(���QP�������ҡt��H�I�U�R������P�ыt��B�P������Q�ҡt��H�A������R�Ћt��Q�J������P�ыt��B�P��x���Q�ҡt��H�A��X���R�Ћt��Q�J��8���P�ыt��B��H���Q�P�ҡt��H�A������R�Ћt��Q�J������P�ыt��B�P��h���Q�ҡt��H�A������R�Ћt��Q�J������P�ыt��B�P��(���Q�ҋE�t��Q��<P���ĉE�P�B�Ћt��Q�E��RP�M�Q�ҋM��������t��H�A��x���R�Ћt��Q�Jj j���x���h�sP�ыt��B�P������Q�ҡt��H�Aj j�������h\tR�Ћt��Q�J������P�ыt��B�Pj j�������h\tQ�ҡt��H�A�����R�Ћt��Q�J��@j j������h�tP�ыV�D:(��j0j �D:�t��H�A$jj ����X����$R�Ћt��Q�J�E�������P�ыt��B�U��@������QR�Ћt��Q�J��X���P����V��,�D:�`�t��H�A$j0j jj ��������$R�Ћt��Q�J�E���8���P�ыt��B�U��@��8���QR�Ћt��Q�J�����P�ыV�t��D:�H�A$��,j0j j�|:j ����8����$R�Ћt��Q�J��������P�ыt��B�P������QW�ҡt��H�A��8���R�Ћt��Q�J�E�P�ыt��B�M�Q������@R�Ћt��Q�B<��8�M��Ћt��Q�RLj�j�������QP�M��ҡt��H�A��(���R�Ћt��Q�R��(���P�M�Q�ҡt��P�B<����(����Ћt��Q�RLj�j�������QP��(����ҡt��H�A��H���R�Ћt��Q�R��H���P��(���Q�ҡt��P�B<����H����Ћt��Q�RLj�j���8���QP��H����ҡt��H�A��H���R�Ћt��Q�R��H���P��H���Q�ҡt��P�B<����H����Ћt��Q�RLj�j�������QP��H����ҡt��H�A������R�Ћt��Q�R������P��H���Q�ҡt��P�B<���������Ћt��Q�RLj�j�������QP�������ҡt��H�A��h���R�Ћt��Q�R��h���P������Q�ҡt��P�B<����h����Ћt��Qj��RLj���x���QP��h����ҡt��H�I�U�R��h���P�ыt��B�P��h���Q�ҡt��H�A������R�Ћt��Q�J��H���P�ыt��B�P��H���Q�ҡt��H�A��(���R�Ћt��Q�J�E�P�ыt��B�P������Q�ҡt��H�A��8���R�Ћt��Q�J������P�ыt��B�P�����Q�ҡt��H�A������R�Ћt��Q�J������P�ыt��B�P��x���Q�ҋE�t��Q��<P�B����W�Ћt��Q�J�E�WP�ыM����C����t��B�P�����Q�ҡt��H�Aj j������h�sR�Ћt��Q�J������P�ыt��B�Pj j�������h\tQ�ҡt��H�A��(���R�Ћt��Q�Jj j���(���h\tP�ыt��B������Q�P�ҡt��H�A��@j j�������h�tR�ЋF�t��Q�J$��j0�|[�j �j��D8�j ����x����$P�ыt��E��B�P������Q�ҡt��H�E��I������RP�ыt��B�P��x���Q����F�d8��,j0j ǡt��H�A$jj ����h����$R�Ћt��Q�J�E���X���P�ыt��B��X���Q�U��@R�Ћt��Q�J��h���P�ыF�t��8��,j0j jǋB�P$j ����H����$Q�ҋ��t��H�A������R�Ћt��Q�J������PW�ыt��B�P��H���Q�ҡt��H�A��X���R�Ћt��Q�R��X���P������Q�ҡt��P�B<��8��X����Ћt��Q�RLj�j�������QP��X����ҡt��H�A��x���R�Ћt��Q�R��x���P��X���Q�ҡt��P�B<����x����Ћt��Q�RLj�j���(���QP��x����ҡt��H�A������R�Ћt��Q�R������P��x���Q�ҡt��P�B<���������Ћt��Q�RLj�j���X���QP�������ҡt��H�A������R�Ћt��Q�R������P������Q�ҡt��P�B<���������Ћt��Qj�j�������Q�RLP�������ҡt��H�A��h���R�Ћt��Q�R��h���P������Q�ҡt��P�B<����h����Ћt��Q�RLj�j�������QP��h����ҡt��H�A�����R�Ћt��Q�R�����P��h���Q�ҡt��P�B<��������Ћt��Q�RLj�j������QP������ҡt��H�I�U�R�����P�ыt��B�P�����Q�ҡt��H��h����AR�Ћt��Q�J������P�ыt��B�P������Q�ҡt��H�A��x���R�Ћt��Q�J��X���P�ыt��B�P������Q�ҡt��H�A��X���R�Ћt��Q�J������P�ыt��B�P������Q�ҡt��H�A��(���R�Ћt��Q�J������P�ыt��B�P�����Q�ҋE�t��Q��<P�B����W�Ћt��Q�J�E�WP�ыM����R����V|�E�<���  �t��H�A�U�R�Ћt��Q�Jj j��E�h�sP�ыt��B�P�M�Q�ҡt��H�Aj j��U�h\tR�Ћt��Q�J�E�P�ыt��B�Pj j��M�h\tQ�ҡt��H�A������R�Ћt��Q�J��@j j�������h�tP�ыF�t���j0�|[	�j �j��D8ǋB�P$j ����(����$Q�҉E��t��H�A������R�Ћt��Q�M��R������PQ�ҡt��H�A��(���R����F�d8�t��Q�J$��,j0j �jj ��������$P�ыt��E��B�P�����Q�ҡt��H�E��I�����RP�ыt��B�P�����Q�ҋF�8��,j0j ǡt��H�A$jj ���������$R�Ћt��Q�J�������P�ыt��B�P�����QW�ҡt��H�A������R�Ћt��Q�J�E�P�ыt��B�@�M�Q������R�Ћt��Q�B<��8�M��Ћt��Q�RLj�j������QP�M��ҡt��H�A�U�R�Ћt��Q�R�E�P�M�Q�ҡt��P�B<���M��Ћt��Q�RLj�j��M�QP�M��ҡt��H�A������R�Ћt��Q�R������P�M�Q�ҡt��P�B<���������Ћt��Q�RLj�j������QP�������ҡt��H�A������R�Ћt��Q�R������P������Q�ҡt��P�B<���������Ћt��Q�RLj�j��M�QP�������ҡt��H�A�����R�Ћt��Q�R�����P������Q�ҡt��P�B<��������Ћt��Qj�j�������QP������RL�ҡt��H�A��8���R�Ћt��Q�R��8���P�����Q�ҡt��P�B<����8����Ћt��Q�RLj�j��M�QP��8����ҡt��H�I�U�R��8���P�ыt��B�P��8���Q�ҡt��H�A�����R�Ћt��Q�J������P�ыt��B�P������Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P�����Q�ҡt��H�A�����R�Ћt��Q�J������P�ыt��B�P������Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҋE�t��Q��<P�B����W�Ћt��Q�J�E�WP�ыM��������E�V|�@;E�E�j����}��t��H�A�U�R�Ћt��Q�Jj j��E�h�tP�ыt��B�P�M�Q�ҡt��H�Aj j��U�hPtR�Ћt��v,�Q�J(������VP�ыt����B�P�M�Q�ҡt��H�A�U�RV�Ћt��Q�J������P�ыt��B�P�M؃�@Q�ҡt��H�I�U�R�E�P�ыt��B�P<���M��ҋt��Q�RLj�j��M�QP�M��ҡt��H�A�U�R�Ћt��Q�R�E�P�M�Q�ҡt��P�B<���M��Ћt��Q�RLj�j��M�QP�M��ҡt��H�I�U�R�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћ]��S����t��Q�BV�Ћt��Q�J�E�VP�у�������S�������t��B�P�M�Q�҃�_^[��]� �������������U���  �t��USVWj ��HH��p  h�  R�Ћt��Q�}��j �E����   j���Ћt��Qj �E����   j���Ћt��Q�J���E�P�}��у�����  �~ ��  ��h�����  �����R�ʛ ���� P��h������  ��������  �t��H�A�U�R�Ћt��Q�Jj j��E�h�tP�у��U�R��h����>�  �t��H�A�U�R�Ћt��Q�J�E�P�ыt��B�Pj j��M�h�sQ�ҡt��H�A�U�R�Ћt��Q�Jj j��E�h�tP�у�,�U�R�E�P�����Q��h������  �����  P�U�R�E�P��?  ��P�M�Q�?  �t��J�U�RP�A�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ѓ� �������  �t��Q�J�E�P�ыt��B�P�M�Q�ҋ]�t��H�Q��S����W�ҡt��H�A�U�WR�Ѓ��������S��������h����"�  ��]�t��Q�J�E�P�ыt��B�Pj j��M�h�sQ�ҡt��H�A�U�R�Ћt��Q�Jj j��E�h�tP�ыt����   �M�Px��(�ҍM�QP�U�R�E�P�k>  ��P�M�Q�^>  �t��J�U�RP�A�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�у�$�t��B�HS����W�ыt��B�P�M�WQ�҃�������S���W����E�}PWS���w����}� t�M��UQRWS���P����t��H�A�U�R�Ћt��Q�Jj j��E�h�tP�ыt��B�P�M�Q�ҡt��H�Aj j��U�h`tR�ЋU��(�M�QR�E�P�t���P�M�Q�U�R�&=  ��P�E�P�=  �t��Q�R�M�QP�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��J�Q��(S����P�E�ҡt��H�U�IR�E�P�у����d����t��B�P��X���Q�E    �ҡt��H�Aj j���X���h�rR�Ћt��Q�J�E�P�ыt��B�Pj j��M�h�rQ�҃�(�} �E    �U  �}� ��  �~ ��  ���   �M�������   �t���� ���   �ȋBx�Ћt��Q�R�M�QP�ҡt��P�Rx����X���P�M��҅��8  �t��H�A�U�R�Ћt��Q�Jj j��E�h�sP�ыt��B�P�M�Q�ҡt��H�Aj j��U�h�tR�Ѓ�(�M�Q�U�R�E�P������Q�;  ��P������R�;  �t��Q�R�M�QP�ҡt��H�A������R�Ћt��Q�J������P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ѓ�$S���ĉE�t��QP�B�Ћt��Q�E�RP�M�Q�҃����W����t��H�I��X���R�E�P�у��t��B�P��H���Q�ҡt��H�Aj j���H���h�tR�Ћt��Q�R�E�P��H���Q�ҡt��H�A��H���R�ЋO|�U�� �<� �E    �o  �]�ۡt��H�A��8���R�Ћt��Q�Jj j���8���h\tP�ыt��B�P<���M��ҋt��Q�RLj�j���8���QP�M��ҡt��H�A��8���R�ЋG4��VÍD�t��Q�J(P�����P�ыt��E�B�P��(���Q�ҡt��H�E�I��(���RP�ыt��B�P�����Q�ҡt��P�B<���M��Ћt��Qj�j���(����RLQP�M��ҡt��H�A��(���R�Ѓ��}� �  �\ �  �t��Q�J�E�P�ыt��B�Pj j��M�h�tQ�ҡt��P�B<���M��Ћt��Q�RLj�j��M�QP�M��ҡt��H�A�U�R�ЋGL��NÍD�t��Q�J(P��t���P�ыt��E�B�P�M�Q�ҡt��H�E�I�U�RP�ыt��B�P��t���Q�ҡt��P�B<���M��Ћt��Qj�j��M��RLQP�M��ҡt��H�A�U�R�Ѓ��E�O|�U@��;��E������]�t��H�A�U�R�Ћt��Q�Jj j��E�h�sP�ыt��B�P<���M��ҋt��Q�RLj�j��M�QP�M��ҡt��H�A�U�R�Ћt��Q��S���ĉEP�B�Ћt��Q�E�RP�M�Q�҃��������E�O|��U@;E�E������t��H�A�U�R�Ћt��Q�Jj j��E�h�tP�ыt��B�P�M�Q�ҡt��H�Aj j��U�hPtR�Ћt��Q�E�R(P��t���Q�ҋ��t��H�A�U�R�Ћt��Q�J�E�PW�ыt��B�P��t���Q�ҡt��H�A�U���@R�Ћt��Q�R�E�P�M�Q�ҡt��P�B<���M��Ћt��Q�RLj�j��M�QP�M��ҡt��H�A�U�R�Ћt��Q�R�E�P�M�Q�ҡt��P�B<���M��Ћt��Q�RLj�j��M�QP�M��ҡt��H�I�U�R�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt���S�����Q�BW�Ћt��Q�J�E�WP�у�������S���4����t��B�P�M�Q�ҡt��H�A��X���R�Ћt��Q�J�E�P�у�_^[��]� U��t���   SV��H�A�U�WR�Ћt��Q�Jj j��E�h\tP�ыt��B�P�M�Q�ҡt��H�I�U�R�EP�ыt��B�P<�� �M��ҋt��Q�RLj�j��M�QP�M��ҡt��H�A�U�R�ЋM�]��QS�U�R���
����t��H�A�U�R�Ћt��Q�Jj j��E�h�sP�ыt��B�P�M�Q�ҡt��H�Aj j��U�h\tR�Ћt��Q�J�E�P�ыt��B�Pj j��M�h\tQ���E���<�E�Pj0j jj ���M��$Q�����E���P�U�Rj0j jj ����x����$P�����E���P�M�Qj0j jj ����\����$R�Z�����P�� ���P�2  ��P�� ���Q�2  ��P��@���R�2  ��P�����P�z2  ��P��0���Q�j2  �t����B�P<���M��ҋt��Qj�j�WP�BL�M��Ћt��Q�J��0���P�ыt��B�P�����Q�ҡt��H�A��@���R�Ћt��Q�J�� ���P�ыt��B�P�� ���Q�ҡt��H�A��\���R�Ћt��Q�J��x���P�ыt��B�P�M�Q�ҡt��H�UЋAR�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҋE�t��Q��,P�B����W�Ћt��Q�J�E�WP�у��������Uh�  RS���<������4  h�  P��P���P���0����M��8�  �M�Q��l����)�  �MP��P���R�E�P��} P�� ���M����  ��l������  �t��Q�J�E�P�ыt��B�Pj j��M�h\tQ�ҡt��H�A�U�R�Ћt��Q�Jj j��E�h�tP�у�(�U�R�EP�M�Q��x���R�E0  ��P�E�P�80  �t��Q�R�M�QP�ҡt��H�U��AR�Ћt��Q�J��x���P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыt��B�Pj j��M�h�sQ�҃�8�E�P��x���Q�M���  P�U�R�/  ���t��P�B<���M��Ћt��Qj�j�WP�BL�M��Ћt��Q�J�E�P�ыt��B�P��x���Q�ҡt��H�A�U�R�ЋM�t��B��Q�H����W�ыt��B�P�M�WQ�҃���������M���  ��P�����  �t��H�A�U�R�Ћt��Q�J�EP�у�_^[��]�$ �U����   SV��W�M����  �t��H�A�U�R�Ѓ��M�Q�Mj�U�R����P��8�����  ��8���P�M��y�  ��8����~�  �t��Q�J�E�P�ыt��B�P�M�Q�ҋM���E�P�Kz P�M��R�  �M��:�  �t��Q�J�E�P�ыt��B�P3�Sj��M�h�tQ�҃��E�P�M���  �t��Q�J�E�P�у��U�R�M���  P膗 �t��H�A�U�R�Ѓ���  h1D4ChCD4C�E����)� PSj�M�Q����  ��u"�U�R�m�  ���M��]���  3�_^[��]� �F;É]�  �F�M�t��<��B�P�M�Q�ҡt��H�A��t���R�Ћt��Q�Jj j���t���h�sP�ыt��B�P��T���Q�ҡt��H�Aj j���T���huR�Ћt����   �Bx��,���Ћt��Q�J�؍E�P�ыt��B�@�M�Q��T���R�Ћt��Q�B<���M��Ћt��Qj�j�SP�BL�M��Ћt��Q�J�E�P�ыt��B�@�M�Q�U�R�Ћt��Q�B<���M��Ћt��Q�RLj�j���t���QP�M��ҡt��H�I�U�R�E�P�ыt��B�P�M�Q�ҡt��H�A�U�R�Ћt��Q�J��T���P�ыt��B�P��t���Q�ҋE��t��Q��P�B����S�Ћt��Q�J�E�SP�у����F����t��B�P��d���Q�ҡt��H�Aj j���d���h�tR�Ћt��Q�R�E�P��d���Q�ҡt��H�A��d���R�ЋM��t��B�� Q�H����S�ыt��B�P�M�SQ�҃���诽��h�  W��袺����tG�t��H�Q����S�ҡt��H�Qj j�h�tS�ҋE��M��h4  h@  WPQ������h�  W���J�����tI�t��B�H����S�ыt��B�Hj j�h�tS�ыU��E��h�	  hD  WRP�������t��Q�J��D���P�ыt��B�Pj j���D���h�tQ�ҡt��H�I�U�R��D���P�ыt��B�P��D���Q�ҋE��t��Q�� P�B����W�Ћt��Q�J�E�WP�у����e����t��B�P�M�Q�ҡt��H�Aj j��U�h�tR�Ћt��Q�R�E�P�M�Q�ҡt��H�A�U�R�ЋM��� Q�t��B�H����W�ыt��B�P�M�WQ�҃����ڻ���t��H�A�U�R�Ћt��Q�Jj j��E�h�tP�ыt��B�@�M�Q�U�R�Ћt��Q�J�E�P�ыU��t��H�� R�Q����W�ҡt��H�A�U�WR�Ѓ����P����M�Q�������t��B�P�M�Q�ҋE@��;F�E������M���  �E�P�/�  ���M��E�    �=�  _^�   [��]� ���������������U���  SVW��hG  �������b� �K 3����������;���  ���������  �t��H�A�U�R�Ћu���M�Qj�U�R�������P�M��.�  �E�P��������  �M���  �t��Q�J�E�P�ыt��B�P�M�Q�ҋM���E�P�ds P�������h�  �M��P�  �t��Q�J�� ���P�ыt��B�PWj��� ���hpvQ�҃��� ���P��������  �t��Q�J�� ���P�у���l������  �t��B�M�Q�P�҃��E�Pj�M�Q��� ���P�M��7�  �U�R��l�����  �M���  �t��H�A�U�R�Ћt��Q�J�E�P�у�hdv�M���  �U�R��l����n�  �M��V�  �������[�  �t��H�A�U�R�Ѓ��M�Qj�U�R���f���P�M���  �E�P���������  �M���  �t��Q�J�E�P�ыt��B�P�M�Q�҃�hXv�M���  �E�P���������  �M���  �M�Q�������l�  P�V� �t��B�P�M�Q�҃��E�P��l����B�  P�,� �t��Q�J�E�P�у��U�R��������  P�� �t��H�A�U�R�����U����U��M��PvQ�]��U�R��x����U�P�荍�����U�Qݝx����������U�ݕ����ݕ����ݕ����ݕ����ݝ����譯���t����   ���   �ыMWP�E��m �t����   �M􋐐   �҅��!  �h�  h1D4ChCD4C�E��E��� �M�PWj������P��  ��uV�M�Q�C�  �t��}����   ���   �M�Q�҃��}􍍈����7�  ��l����,�  �������!�  3�_^[��]� Wh�s�M������E�P�����M�Q�U�R��������  PW�#  ����蛶���t��H�A�U�R�Ћt��Q�J�E�P�у�j h�s�M�覜���U�R�����E�P�M�Q��l����J�  PW�S#  �����9����t��B�P�M�Q�ҡt��H�A�U�R�Ѓ�j h�s�M��D����t��Q���   �}�j j����W�����M�QP�U�R��褷��PW��"  �����õ���t��H�A�U�R�Ћt��Q�J�E�P�ыt��B���   ��3�Wj����;�t�E�P����Wh@v譛�����f����t��Q���   Wj����;�t�M�Q����Wh0v�x������1����t��B���   Wj����P�E�P���߶��P��� �t��Q�J�E�P�ыM����\�  Wh v�M�����Whv�M������U�R�����P��������  P�M�Q������R�!  ��P������P�!  P胋 �t��Q�J������P�ыt��B�P������Q�ҡt��H�A�����R�Ћt��Q�J�E�P�ыt��B�P�M�Q�҃�$�9�  h1D4ChCD4C�E��E��ԉ �M�PWj������P�Q�  ��u(�M�Q��  �U�R�}���  ���M�}��J  ������t��H�A�� ���R�Ѓ�Wh�u�M������t��Q�R�� ���P�M�Q�ҡt��H�A�U�R�ЋM���Q���� �����R�~������g����   �E��E��E�P�E��  �}��}��}��� ��Wh�s�M��r���Wh�u�M��d����M�Q�U�R�����h�uP��� P�M�Q������R�
   ��P������P��  ��P�� ���������t��Q������P�J�ыt��B�P������Q�ҡt��H�A�����R�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҋE���P���� �����R�q������Z���Wh�s�M�茘��Wh�u�M��~����t�� �M�QP�����R�v���P�E�P������Q�%  ��P������R�  ��P�� ��������t��H�A������R�Ћt��Q�J������P�ыt��B�P�����Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�ыU���R���� �����P荗�����v����M�Q�������t��B���   Wj���ҋM�{�{�Eȡt����   ���   �}��Ѕ��e  ��� �t����   �E��M􋒔   P�ҋ��t����   �B�ω}���=�  ��  �t��Q�J������P�ыt��B�Pj j�������h�uQ�ҡt����   �Bx������P������Q������R�  P臈 �t��H�A������R�Ћt��Q�J������P�у������������t��B�P������Q�ҡt��H�Aj j�������h�uR�Ћt����   �Bx������P������Q������R�  P�ކ �t��H�A������R�Ћt��Q�J������P�у��}� ��  �t��BH���   h�  ��V�у�P��<����   j��T�����  j ��<����  ���E�    �� ���}�����  �	��$    ���t����   �P����=�  �|  hF  h�  W���P������b  j ���E�   �H� ������  h�  W�E�P��������t��Q�B<�M��Ѕ���   V��T����x  �M���� ������   ��    �t����   �B����=)  ��   �t����   �Bx���Ћt��Q�Rx�M�Q���҅�ue���и �M�Q������R3�V�ȉE��� ��tB�d$ ������F;E��d$ ��h�����@���I��@;E�~�E�P������Q�M�V�V� ��ut����   �P(���ҋ����5������X���j ��<����0�n  �t��Q�J�E�P�ы}����t����   �P(���ҋ��E����F�����X����8 ��   �t��Q�J�E�P�ыt��B�Pj j��M�h�uQ�ҡt����   ��������R|���E�P�ҡt��H�A�U�R�Ћ�t��QT3�WP�B�Ѓ�;���  �����Q���}� ��t��U��U��M��]�Q�B�PHh�  ������ҋ�X�������������  �}� ��   ��h��� �E�    ��   ��3�9s~]���$    �S�t���� ���   �ȋBx�Ћ�X����U������t����   �Bx�Ћt��Q�ȋBxW�Ѕ�t1F;s|��s��X����U��<���|jjjV����  ��t�C�<��E�@;�h����E��^����t��QH�u܋�p  j h�  V�Ћt��QHj �Eċ�p  h�  V�Ћt��QH���������   h�  V�Ћt��QH�����   h�  V�}��Ћ���4�����(�u�;�t(}+�PV�� ����:  �jj��+�QP�� ����#  3���~;���������d$ �������3�;Q��$�����@����;Ɖ\��������|Ջ}�������P���t�����8���������;�t ������}+�PW�  �jj+�WP�  �t��QH�M܋R8��X���P�ҋ�   �����������P������Q��$���R�s�����݅|���3ۃ}�݅t���݅l���݅d���݅\���݅T����  �}��Uă���B(����G��    ݅<����������H؍t��܅$������H������H����]�݅D����H�܅,������H������H����]�݅L����H�܅4������H������H����E���E��Y�Y������݅<����L1�H�܅$������H���������]�݅D����H�܅,������H���������]�݅L����H�܅4������H���������E���E��Y�Y݅<����H܅$������H�����H���������L��]�݅D����H܅,������H�����H���]�݅L����H܅4������H�����H���E���E��Y�Y������݅<����L �H ȃ�`��܅$������H������H���ݝ����݅D����H�܅,������H������H���ݝ���݅L����H�܅4������H������H���݅�����]�݅������]��E���Y�E��Y����;]���   �Mč[�D��U�����+�+�݅<����������H��ȃ���܅$������H������H���ݝ����݅D����H�܅,������H������H���ݝ���݅L����H�܅4������H������H���݅�����]�݅������]��E���Y�E��Y�e�����8����݋���������������;�t&}+�QP�������3  �jj+�PQ�������  �]�3�3Ʌ�~}��������$������d$ �<�������u.�r�4��2�������t��r��������t��r��������t���2�4��r��������t��r��������t���$����A��;�|��t��B�M���   j j�҅��X  �t��HH�u܋��   j h'  V�ҋ������[  ��8���������;�t,}+�QP�������-  �jj+�PQ�������(  ��8��������;�t&}+�QP��������	  �jj+�PQ��������  ���˷ ��ݕ$���3�ݕ,���3�ݕ4���������ݕ<���ݕD���ݕL���ݕT���ݕ\���ݕd���ݕl���ݕt���ݝ|������a  �t��HD�������I,��$���RWP�ы�$����v�Ƀ�Ƀ<��7  ��������l������p����T��t����T��x����T��|����T�U��T��������D��T������X����P��\����H��`����P��d����H��h����P�������N�I��<������@����P��D����P��H����P��L����P��P����P�������V�R�Ë�$������(����X��,����X��0����X��4����X��8����X�������4��������F�D��������]�������������   �������
��T������X����P��\����P��`����P��d����P��h����P�������D��<������@����P��D����H��H����P��L����H��P����P�������N�I��$������(����P��,����P��0����P��4����P��8����P�������4��������V�T�����������$���4�G;�������M��E��}������SQ�M܍�����RPQW�������������V�t��P���   j j���Ѕ�t	������N������販���ދ��t��}����   �M􋐐   G�}���;������3��M��.�  9}�t9{~�EVP�������t��Q�J�� ���P�эU�R��  �E�P�}���  ���  j h�u������褈��3�Vh|u�M�蔈���t����   �M܋Bx�Ѝ�����QP�U�R������P�9  ��P������Q�)  P�y �t��B�P������Q�ҡt��H�A������R�Ћt��Q�J�E�P�ыt��B�P������Q�҃� �������u����t��H�A�� ���R�ЍM�Q��  �U�R�u���  ���M�u���  �w����������.����t��H�A�� ���R�ЍM�Q�q�  �U�R�}��e�  �t��}����   ���   �U�R�Ѓ������t��Q�J�E�P�ыt��B�P3�Wj��M�hHuQ�ҡt��H�A�U�R�Ћt��Q�JWj��E�h<uP�ыt����   �Px��(���ҋ�t��H�A������R�Ћt��Q�R������P�M�Q�ҡt��P�B<���������Ћt��Qj�j�VP�BL�������Ћt��Q�J�����P�ыt��B�@�����Q������R�Ћt��Q�B<��������Ћt��Q�RLj�j��M�QP������ҍ����P��v �t��Q�J�����P�ыt��B�P������Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�у��������I����t��B�P�� ���Q�ҍE�P��  �M�Q�}���  �t��}����   ���   �M�Q�҃��7����t��Q�J�E�P�ыt��B�PWj��M�h$uQ�ҍE�P��u �t��Q�J�E�P�у�������R薨 �t����   ���   �U�R�Ѓ��������}����  ��l�����  ��������  _^�   [��]� ���������̡t�V�񋈈   ���   V�҃��    ^���������������U��Q3�9A~V�u�2@��;A|�^]� ���������������U��EV���
�   ^]� �MW��|/�~;�}(�> t#�~ u%�t��H��0  h�sh�  �҃�_3�^]� ��;�|���k���_�   ^]� S�;�|�ߋ�+���;ȉ]��   ^��~�F�I���QP�[��P��` ���N��~;ύI�ЉV�'  ������V+ӍR���R��)F+ȍ@��N�N�Q�+�Q�` �F�t��Q���  �@�h�s�h�  �PQ�҃������   �N)^�I[��_�V�   ^]� �V��+Ë^�D�����W�@��;ʋ]�E}-�F+�+�����R��R��R�I��R��_ �E��;F}L�t��Q���  �@�h�s�h�  �PQ�҃����u	[_3�^]� �N�I�ȋE�F�V)^[_�   ^]� ��U��EV���
�   ^]� W�}��|/�N;�}(�> t#�~ u%�t��H��0  h�sh�  �҃�_3�^]� ��;�|���k���_�   ^]� S�;�|�ً�+���;��]��   ^��~�F��    QP��R��^ ���N��~;ύ��V��   ������V+���R��)F+ȉN�N�Q�+�Q�^ �F�t��Q���  h�s�h�  �PQ�҃������   �N)^[��_�V�   ^]� �V��+ÍD���~��C�^�A�;�}!�U�F+�+���Q׍�Q��R� ^ ��;^}C�t��H���  h�sh�  ��    RP�у����u	[_3�^]� �V���F�^�])^[_�   ^]� ���U��t��P�B<V���Ћt��Q�M�RLj�j�QP���ҋ�^]� �������������U���VW�}���}
_3�^��]� S�]����  �F;ǋ��ύ�N�U��u(�t��H��0  h�shA  �҃�[_3�^��]� ��;���  )^�F�Y  @���j j�и   +�����؋F�ʙÉ]����SP�E��C` �ȉU��;�u��E�;�u�;�|�;M�r��]�Ù9U�E�|�;��{����F�U��NF�@����N��h�s��u�t��Q���  hW  P�у���t��RhX  PQ��  �у��ȉ�������F�@�F�щN��~N+Ǎ@���P��+E�Í@��P��@��P��[ +]��F����Q�[��QP��[ ���}  �@�ҋ�+E��R�@���[R��Q�[ ���V  ��~�N����R�@�Q��Q�[ ���F�@��ЉN�   �F�D����@����؋F�ʙ;ʉM���   ;���   j jQS�^ �ȉU��;������E�;�� ���;E������;�������E�9U�E������;�������h�s��u%�t��Q���  �[���h|  P�у��$�t��J�[��h}  �RP��  �Ѓ��ȉ���s����F�@�щF�^�F;�}*�N+Ǎ@���R����E�R�@��P�ZZ ���]�} tG�N;�}"��+��@���R�I�N��j R�(Y ���V�[���P���j P�
Y ���} tO�N��;�}!�F�I�Ћ�+х�t��P�P����u�V��ʅ�~�˅�t��P�P����u��؋E�F[_�   ^��]� ��������������U���VW�}���}
_3�^��]� S�]���  �F;ǋ��ύ�N�U���u(�t��H��0  h�shA  �҃�[_3�^��]� ��;��h  )^�F�.  @���j j�и   +�������F�ʙ��߉}���WS�T\ �ȉU�;�u��E�;�u�;�|�;�r��]�Ù9U�|�;�r��M�F�V��Fы���Vh�s��u�t��Q���  hW  P�у���t��RhX  PQ��  �у�����!����V�}�N���F��~>+�ɋ�+U��QӍ��Q��P�$X �F+]��    Q��RP�X ���V  �ɋ�+U�Q��Q��R��W ���7  ��~�V��    Q�R��R��W ���F����V�	  �F�D����@����؋F���;���   ;���   j jWS��Z �ȉU�;��A����E�;��6���;��.���;��$����E�9U�����;������h�s��u#�t��Q���  ��    h|  P�у��"�t��Jh}  ��    RP��  �Ѓ����������N���V�^�F9E}"�M�V+���P��P�Eȍ�Q�V ���}�} t=�F;�}�N��+���R��j R�U ���E�V��    Q��j P�nU ���M��N[_�   ^��]� �������U��t��H�QV�uV�ҡt��H�U�AVR�Ћt��Q�B<�����Ћt��Q�M�RLj�j�QP���ҋ�^]���������U��Q�E;�u	�   ]� }+�RP�?���]� jj+�PR�.���]� ����������U��V��W�~��}_3�^]� jjjW�������t�F�M��_�   ^]� �������xv��Y �����U��V���xv�Y �Et	V�C? ����^]� ���������U��M�UV�uW��r�;u��������s��tE��9+�u1��v6�B�y+�u ��v%�B�y+�u��v�B�I+���_��^]�_3�^]�����������U��QV��j �M��GG �F���s@�F�M��[G ^��]�������U��QVW��j �M��G �G��v	���sH�G�w����֍M�#��G _��^��]������v����������U��QW�9��t=j �M���F �G��v	���sH�GV�w����֍M�#���F ��t
��j����^_��]����U���EV����vt	V��= ����^]� �������������̰�������������̸   �����������U��A$V�0W�}j �M�7�F �F���s@�F�M�3F ��_^]� �����������U��MV3��� ��t�t����   ���ȋB(�Ѕ�u��^]� ��������������U���SVW���� �O ���EP�2F P���� �M��B�  �t��Q@�J$�E�PV�ыt��B�P4��jh�  �M��ҡt��P�B4jh�  �M��Ћt��E�Q�R8Ph�  �M��ҡt��P�B4jh�  �M��Ћt��Q@�J(j�E�PV�ы]����3��� ��t�d$ �t����   ���ȋB(�Ѕ�u�WV���~� �t����   �Bj j���ЍM���  �t��Q�J�EP�у�_^[��]� �U���4�t��UV��HT�Aj R�u��Ѓ��E��u^��]� S�M�Q���ġ ���   +��   �]�ƨ   ���Q���������;�r�|Y �t��Q�F�RHW��i��   �L8 Qh�  �M��ҋN+N���Q���������;�r�5Y �N��9�    _tSS����M  �t��R��P�B8h�  �M��ЋM���Q�M��O�  �t��B�P<�M�Qh�  �M��ҍM�譮  �M�E�P�� �M��y�  [�   ^��]� ������������U���L�t�SVW���H�A�U�R�}��Ћt��Q�Jj j��E�h�rP�ы��   +��   �]�Ǩ   ���Q���������;�r�;X �t��Q�Rx��i��   G�M�Q���   �ҋ�t��H�A�ލU��R���Ѓ����v  �t��QT�u�Bj	V��3Ƀ��E;�u_^3�[��]� Q�M�M�M�Qh�  �M�誉 P���� �M��J{ �t����   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   �^� P���� �M���z �t����   �
�E�P�у��u�U�R���I� S���L  �t��Q��PP�BHh�  �M���S����K  ���    tUS����K  �t��Q�   P�B8h�  �M��ЋM���Q�M��#�  �t��B�P<�M�Qh�  �M��ҍM�聬  �E�P���� �M��N�  �t����   �
�E�P�у�_^�   [��]� ���������U���L�t�SVW���H�A�U�R�}��Ћt��Q�Jj j��E�h�rP�ы��   +��   �]�Ǩ   ���Q���������;�r��U �t��Q�Rx��i��   G�M�Q���   �ҋ�t��H�A�ލU��R���Ѓ����T  �t��QT�u�BjV��3Ƀ��E;�u_^3�[��]� Q�M�M�M�Qh�  �M��j� P���Ҏ �M��
y �t����   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   �� P��覎 �M��x �t����   �
�E�P�у��u�U�R���	� S����I  ���    tUS���I  �t��Q�   P�B8h�  �M��ЋM���Q�M���  �t��B�P<�M�Qh�  �M��ҍM��c�  �E�P���Ȝ �M��0�  �t����   �
�E�P�у�_^�   [��]� �����������U���L�t�SVW���H�A�U�R�}��Ћt��Q�Jj j��E�h�rP�ы��   +��   �]�Ǩ   ���Q���������;�r��S �t��Q�Rx��i��   G�M�Q���   �ҋ�t��H�A�ލU��R���Ѓ�����  �t��QT�u�BjV��3Ƀ��E;�u_^3�[��]� Q�M�M�M�Qh�  �M��J� P��貌 �M���v �t����   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   ��� P��膌 �M��v �t����   �
�E�P�у��M�U�R�� S���G  ـ�   �5�vj �E�Ph  �M��E�   �]�E�]�蔄 P���� �M��4v �t����   �
�E�P�у�S���EG  ���    tUS���4G  �t��R�   P�B8h�  �M��ЋM���Q�M�艧  �t��B�P<�M�Qh�  �M��ҍM���  �M�E�P�K� �M���  �t����   �
�E�P�у�_^�   [��]� ��������������U���L�t�SVW���H�A�U�R�}��Ћt��Q�Jj j��E�h�rP�ы��   +��   �]�Ǩ   ���Q���������;�r�[Q �t��Q�Rx��i��   G�M�Q���   �ҋ�t��H�A�ލU��R���Ѓ����T  �t��QT�u�BjV��3Ƀ��E;�u_^3�[��]� Q�M�M�M�Qh�  �M��ʂ P���2� �M��jt �t����   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   �~� P���� �M��t �t����   �
�E�P�у��u�U�R���i� S���!E  ���    tUS���E  �t��Q�   P�B8h�  �M��ЋM���Q�M��e�  �t��B�P<�M�Qh�  �M��ҍM��å  �E�P���(� �M���  �t����   �
�E�P�у�_^�   [��]� �����������U���  ��3ŉE�SVW���CL ��ݕ������`���ݕ�����������PvPݝ����������Q������ݕ����R�荅����ݕ����3�ݝ����P��������l���ݕ����ݕ����ݕ����ݕ����ݕ ���ݝ����{���t��Q�J��L���P�ыt��B�PVj���L���h�wQ�ҍ�L���P�^[ �t��Q�J��L���P�ы��   +��   �����������������h����B
  ��d������   +��   ���������������9�h���r�PN ���   �d����{ �   �}��t{�t��B�P������Q�ҡt��H�Ij j��U�R������P�ы�`�����������R�G9 ��\����t��H�A������R�Ѓ���\��� t��\���Q�5� ���U�E�RP腯 ������x������~	  ���   +��   ���������������9�h���r�mM �t��B���   �P�d���������Q�ҡt��H�Aj j�������WR�Ћt����   �R|��������P���ҡt��H�A������R�Ћt��QH���   j h�  V�Ћt��QHj �E����   h�  V�Ѓ��}� ǅ|���    ~d3ɐ�U�t��l���+���p����t+���t����t�+׉��t���+��p�P��p����P��|���B�� ��;U艕|���|���x���3�9}���   ��l���݅���݅(����M�݅ ����R݅�����ҋ��   ݅������G��܅�������@܍ ��������H��݅�����܅�����@܍��������H��݅�����܅�����@�������H�����Y��Y��Y�;}�|��������؃; �P  �}� �F  ��E�ݕ0���Pݕ8���ݕ@���ݕH���ݕP���ݕX���ݕ`���ݕh���ݕp���ݕx���ݕ����ݝ������� ��3҃���t���;��  9U艕p�����   ��|����
�d$ ��|����M�t
���   �4v�4�V�t
�4v�4�V�t
�L
�4v�I�4���VR��p����jw����   ��0���󥋍t���� � �t��QD��p����R0��0���QVP�҃�|��� F��;u艵p����i�����t�����x���j W��賘 �t����   �Bj j����j h�  ���?� ����   �t��Q�J�� ���P�ыt��B�Pj j��� ���h�wQ�ҡt����   �Bx�����Ћt��Q�J����,���P�ыt��B�@��,���Q�� ���R�Ћt��Q�B<����,����Ћt��Qj�j�WP�BL��,����Ѝ�,���Q��T �t��B�P��,���Q�ҡt��H�A�� ���R�Ѓ��{ �>  �t��Q�J��<���P�ыt��B�Pj j���<���h�rQ�ҋ��   +��   ���Q�鋋�   +��   ������������QuZ���������u��H ���   �t���<���P���U��Q�B��W�Ћt��Q�E��JWP�у�V���k����c  ����������N  ���   +��   ���Q���������u�DH ���   �t���<���P���U��Q�B��W�Ћt��Q�E��JWP�у�V����������   +��   ���Q���������   �;���  ǅ|����   h)  草 �t��Q������t������~  �J������P�ыt��B�Pj j�������htwQ�ҡt��H�A(������WR�Ћt��Q�J�E�������P�ыt��B�U��@������QR�Ћt��Q�J������P�ыt��B�P��L���Q�ҡt��H�I��L���R������P�ыt��B�P<��8��L����ҋt��Q�RLj�j�������QP��L����ҡt��H�I��<���R��L���P�ыt��B�P��L���Q�ҡt��H�A������R�Ћt��Q�J������P�ыt����   �P|����<���Q���ҋ��H� 3�9u�E�~�E�9<�u	�M�V�M� F;u�|鋍x���3��ʔ ��t��    �t����   ���ȋB(�Ѕ�u狍x���V��t���V�4� �t����   �Bj j���Ћ��   +��   ���Q���������;�r�E �t����   �|�����<���R�Q���ĉE�P�B�Ћt��E��Q�JPV�ы�x�����R���9������   +��   ��|����   ���Q��������G�;��R�����x����t��Q�J��<���P�у���`���j j j V���W- �t����   �Pj j����3������������� �����(�����$��������Ph�   ������������Q ������   �M��l���������Tf ���   +��   ��h�����d���x��������������F�h���;�������   _^[�M�3��; ��]ËJ��<���P�у�3�_^[�M�3���: ��]Í������e �M�_^3�3�[��: ��]����U���SV�񋎸   +��   ���Q��������3��W�'  �]����   +��   ���Q���������;�r�C ���   E��N P�. ����ughG  襁 ��������   ���   +��   ���Q���������;�r�9C �t����   ���   E��R|P���ҋN j j W�H+ WS������WS���V����~ W��Su���������WS������jj���\� �t����   �Bj j���Ћ��   +��   �E��   ���Q��������C�;������_^�   [��]Ët��B�P�M�Q�ҡt��H�Aj j��U�h�wR�ЍM�Q��M �t��B�P�M�Q�҃�_^3�[��]�����������V�񋆈   WP�P$ ���   Q�D$ ���   �����n  �R��# ���   3���;�t	P��# �����   P���   ���   ���   �# ���N\苗  �N@胗  �N$�{�  �t��Q�B��V�Ѓ�_^����U��t���S�ًH�AV�SWR�Ѓ��K$�I�  �K@�A�  �K\�9�  j���   �<! 3Ƀ�;�t�0�3�j��N�N�N���   �! 3Ƀ�;�t�8�3���O�O�O�Kx�K|���   ǃ�   �����F�E�9Fv��@ ��M��N�M�;Nv��@ �M��U��R�U�RQP�E�P����_  �w9wv�@ ��M��O�M�;Ov�@ �M��U��VRQP�E�P���}l  _^��[��]�����U���`  ��3ŉE�SV�uW�ٿ   W��X�����  j@WV��`�����  ��u+��X����H��`�����X������y( u��j P�q  ������ �p  �t��Q�J������P�ыt��B�Pj j�������h�xQ�ҡt��H�A��H���R�Ћt��Q�Jj j���H���hvP�ыt��B�P��8���Q�ҡt��H�Aj j���8���VR�Ѓ�<������Q��8���R��H���P��(���Q�������P�����R�����P�J �t��H�A�����R�Ћt��Q�J��(���P�ыt��B�P��8���Q�ҡt��H�A��H���R�Ћt��Q�J������P�у�$��������{  ������Rǅ�����v�O- ��3�_^[�M�3��d5 ��]� �t��H�A������R�Ћt��Q�Jj j�������h�xP�э�����R��J �t��H�A������R�Ћ�X����A����`����c  ���$    �d$ j
��X�����q  ��Rjc������P��X����
�  j������QhXt�M ����uG{|���   +��   ���   ���������������;�r�= ���   ����+΍D�h�  j������Ph�x�-M ����uJ��   ���   +��   ���   ���������������;�r�2= ���   ����+֍D�l�R  j������Qh�t��L �����  ��   jxP������R��3 ���   ��l�����   �   ������@�P���z  ���   +��   ���   ���������������;�r�< ���   ����+�3��|�d���   +��   ���   ���������������;�r�S< ���   ����+Ή|�h���   +��   ���   ���������������;�r�< ���   ����+Ή|�l�   �4j������Ph�x�K ����u���   {xQ���   �f0  ��d8��X����B��`����������`����h  ��u+��X����H��`�����X������y( u��j P�m  �s|3ɋƺ   �������Q�U �����t�V���|�H�Q������Q��Q�y��3����   �؉��   3ɋƺ   �������Q� 3���;�t!�V�;�|��H�Q������Q��Q�y����3����   ���   +��   ��������������3���C  ���   +��   ���������������;�r�: ���   ǋ@d3�@�    �������Q�d ���   +��   ���������������������;�r�:: ���   �������Tp���   +��   ���������������;�r�: ���   ǋ@d3�@�   �������Q�� ���   +��   ���������������������;�r�9 ���   �������Tt���   +��   ��������������F�x;������3���X����QǄX����x������ ǅ`����w��   9�����t��`����Y  ������P�lH ����h�����p�����l�����x�����|�����t����������������`�������������ƅ���� ƅ���� ��������������l�����|�����������h�����x���������������������������������ǅ`����v������;�tU�0;�t@W�������# �F;�v	���sH�F�^����Ӎ�����#��
# ;�t
��j���Ћ�����Q�  ����d����&' ��X����B������ǄX����vQǅ�����v�& �M���_^3͸   [�. ��]� �������������U����  ��3ŉE�SVW��j������k}  ��,����N\P�������&�  �t��Q�Bdj��,����Ћt��Q�����   hzGh�  W�Ћt��Q��j�؋BhWS��,�����j@jS������w  ��u+������I�������������y( u��j P�h  ��X��� �a  �t��B�P������Q�ҡt��H�Aj j�������h�xR�Ћt��Q�J��p���P�ыt��B�Pj j���p���hvQ�҃�(������P��L���Q��������  P��p���R��<���P������P��`���Q�����P��A �t��B�P��`���Q�ҡt��H�A��<���R�Ћt��Q�J��L���P�ыt��B�P��p���Q�ҡt��H�A������R�Ћt��Q�J��,���P�у�(��\�����r  ��\���Rǅ\����v�[$ ��3�_^[�M�3��p, ��]át��H�A��p���R�Ћt��Q�Jj j���p���h zP�ыt��B�P������Q�ҡt��H�Aj j�������h�yR�Ѓ�(��p���Q��������`���R觋  P������P��<���Q������P��L���R����P�m@ �t��H�A��L���R�Ћt��Q�J��<���P�ыt��B�P��`���Q�ҡt��H�A������R�Ћt��Q�J��p���P�у�$������B���������+  �8�����������
��$    �I ������j
�������g  ��Ph�   ������Q������A{  j������Rhu��C �����	  ���   ���   ��������G���   �s)  �GP���r  ������Q������h�yR��D �t��H�A������R�Ћt��Q�Rj j�������P������Q�ҋK+K���Q��������� ;�r�`3 �C�t�������Q�RP������Q�ҡt��H�A������R�ЋK+K���Q��������ʃ�;�r�
3 �S������Ǆ�       �  j������Qh�y�B ����uJ���   +��   ���Q���������;�r�2 ���   �TR������h�yP�C ���A  j������Qh�y�:B ����uJ���   +��   ���Q���������;�r�M2 ���   �TR������h�yP�KC ����  j������Qh�y��A ����uJ���   +��   ���Q���������;�r��1 ���   �TR������h�yP��B ���y  j������Qh�y�rA ����uC���   W���v&  ��0PW���j&  ��(PW���^&  �� P������h�yR�B ���  j������Ph�y�A ����uC���   W���&  ��HPW���&  ��@PW���&  ��8P������h�yQ�-B ���  j������Rh�y�@ ����uC���   W���%  ��`PW���%  ��XPW���%  ��PP������h�yP��A ���b  j������Qh|y�[@ ����uC���   W���_%  ��xPW���S%  ��pPW���G%  ��hP������hlyR�sA ���  j������Phdy��? ����uV������Q������hXyR�9A ��j ������P��`�����J����`���Q���   W����$  �ȃ��^����`����qj������PhPy�? ����u{������Q������hDyR��@ ��j ������P��p����qJ����p���Q���   W���\$  �ȁ��   �/^����p����t��B�PQ�҃�W���/$  ǀ�      ������@����������������3\  ��u+������I�������������y( u��j P�`  j�������t  �������^@R���v�  �t��P�Bdj�������Ћt��Q�����   hzGh  W�Ћt��Q��jW��\���P�Bh�������Ћ�\���j@jQ�������Kn  ��u+�������J���������������y( u��j P��_  ������ �t��H�A��p���R��  �Ћt��Q�Jj j���p���h�xP�ыt��B�P������Q�ҡt��H�Aj j�������hvR�Ѓ�(��p���Q��`���R���S�  P������P��<���Q�O�����P��L���R�?���P�9 �t��H�A��L���R�Ћt��Q�J��<���P�ыt��B�P��`���Q�ҡt��H�A������R�Ћt��Q�J��p���P�ыt��B�P������Q�҃�(�������/j  ��������vP������� �t��Q�J��,���P�у���\�����i  ��\���R��\����q ��3�_^[�M�3��# ��]��Ћt��Q�Jj j���p���h zP�ыt��B�P������Q�ҡt��H�Aj j�������h�yR�Ѓ�(��p���Q��`���R���ӂ  P������P��<���Q�������P��L���R����P�7 �t��H�A��L���R�Ћt��Q�J��<���P�ыt��B�P��`���Q�ҡt��H�A������R�Ћt��Q�J��p���P�ы������B3���$�������������f  j
�������B_  ��Ph�   ������Q�������r  ���   +��   ���Q��������3����   �������t��Q�J������P�ыt��B�@j j�������Q������R�Ћ��   +��   ���Q��������ʃ�;�r��* �t��B���   ������@x������R�Ћt��Q�J���ߍ������PG�у���u2���   +��   �������   ���Q��������C�;��.����������������j������Qh4y� : �����  ���   +��   ���Q���������;�r�* ���   ��i��   ���   R������h$yP�; �������I��j
�������]  ��Rh�   ������P��������p  �t��Q�J��p���P�ыt��B�@j j�������Q��p���R�Ћ��   +��   ���Q��������ʃ�;�r�U) �t����   �B���   R�P��p���Q�ҍ�p�����   j	������Qhy��8 ������   �������Jj
�������\  ��Ph�   ������Q������� p  �t��B�P��`���Q�ҡt��H�Ij j�������R��`���P�ы��   +��   ���Q���������;�r�z( �t��Q���   �R��i��   ���   P��`���Q�ҍ�`����t��H�AR�Ѓ��������A�����������3�������9�����t ����G  ��u3�������R�<7 ����t3��������������������������������������������������`�������������ƅ���� ƅ���� ������������������������������������������������������������������;�u)�������I��������������9y(u��WP��X  ��\���V�7 ������5  �t��B�P��p���Q�ҡt��H�AWj���p���hyR�Ћt��Q�J������P�ыt��B�PWj�������hvQ�ҡt��H�A��`���R�Ћt��Q�JWj���`���VP�у�<��p���R��`���P������Q��<���R������P��L���P�����P��1 �t��Q�J��L���P�ыt��B�P��<���Q�ҡt��H�A��`���R�Ћt��Q�J������P�ыt��B�P��p���Q�҃�$�t��H�A������R�Ѓ���������b  ��������vQ�������b �t��B�P��,���Q�҃���\����b  ��\���P��\����- �M���_^3͸   [�? ��]�������V���������a����   ^�����������U���SVWj�  �]3���;�t��3�jV�M��EQ�M�s�s�s�E�)  �������   �U�U�M��+�PVQ�M��E�   �E�    �E� �Y>  �U�R���u  �}�r�E�P� ��j�wV�MQ�M�:)  �����u��UPVR�M��E�   �E�    �E� �>  �E�P���8u  �}�r�M�Q�I ��_^��[��]� �����������U���X  ��3ŉE�SV�uW��j������������� 3ۃ�;�t��������������������j�������������������� ��;�t��������������������j�������������������������^i  j@jV�������^c  ��u)�������H��������������9Y(u��SP��T  9�0�����  �t��Q�J������P�ыt��B�PSj�������h�xQ�ҡt��H�A������R�Ћt��Q�JSj�������hvP�ыt��B�P������Q�ҡt��H�ASj�������VR�Ѓ�<������Q������R������P��x���Q�A�����P������R�1���P�. �t��H�A������R�Ћt��Q�J��x���P�ыt��B�P������Q�ҡt��H�A������R�Ћt��Q�J������P�у�$��4����6_  ��4���Rǅ4����v� ���������d  �������d  3�_^[�M�3�� ��]� �t��H�A������R�Ћt��Q�JSj�������h zP�ыt��B�P������Q�ҡt��H�ASj�������h�zR�Ћt��Q�J������P�ыt��B�PSj�������VQ�҃�<������P������Q������R������P������P��x���Q����P�, �t��B�P��x���Q�ҡt��H�A������R�Ћt��Q�J������P�ыt��B�P������Q�ҡt��H�A������R�Ћt��Q�J���������P�������������ыt��B�P������Q�������ҡt��H�ASV������h�zR�Ѝ�����Q��, �t��B�P��������@Q�ҋ������@������������	  3����������������$    j
�������S  ��Qh�   ������R��������f  j������Ph�t�k/ ������   ������Q������h�zR�0 ��������P��l����t  ��l����_\Q���kx  ��l����0u  ���w  ������R��l����Wt  ��l���P���x  ��l�����t  �  j������Qh�t��. �����  �t��B�P������Q�ҋ���������������;�v�� ��������������������;�v� ������SVWP������Q��������b  ������ǅ����   ǅ����    ƅp��� �P�@��u�+�P������R��l�����8  jj��l���P��x�����d  ������r��p���Q�(  ��������R�� ���     �@   �@    �� �@ ��x�����P��m  ������Q�p  ������������+˸�$I�����������H��w� �������{4r�[ ��� �t��Q�J������P�ыt��B�Pj j�������SQ�ҡt��H�I������R������P�ыt��B�P������Q�ҋ��������   +��   �ƨ   ���Q���������� 3��tg3ې�N+N���Q���������;�r�� �t��B�N�@x�������R�Ѕ���  �N+N���Q��������Gʁ��   ;�r��N+N���Q�������   ���̍|�&  W���^[  �N+N���Q���������|
��N+N���Q���������;�r�L �t�i��   ~�Q�J������WP�ыN+N���Q���������L���������x����BǄx����w�E��E�wt�M��R���  ���E��     �M��    �U��    �E��     �M��    �U��    �E��e���E�    �E��v����tP���tAj ������� �C��v	���sH�C�s����֍�����#�� ��t
��j����W�7�  ���M��@
 ��x����H�U�Ǆx����vR�EȌv��	 �t��H�A������R�Ѓ��[  �����������j������Qh�t�* ����u9������@P���   �������������H  P������h�zR�+ ���  j������PhXt�B* ����u8���   ��������HQ�PRP������h�zP�l+ ���������  j������Qh�x��) ����ud���   ��HQP������h|zR�$+ ���   ƍHQ�PRP������hlzP�+ �苏�   �d�D��$����������;  j������Rh�x�r) �����  ���������t������P���   �#  �Ht�������4���������^  ������P��l����?  jj��l���Q��x�����_  ��l����9.  ������R�� ���     �@   �@    �� �@ ��x�����P��h  ��h���Q�(k  ��H�������j^  ��������������+˸�$I�����������   �;��>  �����������   �������������j/V�������  P��p���R���M���P�������ac  ��p����Z  j �������y  �xr�@���P�) �x����������Ð   P����  �Hp�������|�j�������1  �Hj h�rQj ���m  ��tJj�������  �xr�@���P�) ��������R�ˍx��d  �������@p���Ή|���������������������+˸�$I����������F�;������+���$I�������������   j �������q  �xr�@���P�( ���������������������ǐ   Q�ύX����  �Pph�rj�������\2�  P�-  ����t<j�������  �xr�@���P�( �X���������P���Y  �Hp�\1�������M���"  �U�R�EȌv�R ��������������3ۋ������@�����������������9�0���t ���76  ��u3���0���Q�% ����t3��������������������������� ��������������������`�����������ƅ,��� ƅ%��� ������������������ ���������������������������0�����(����� ���;�u)�������H��������������9Y(u��SP�G  �t��Q�J������P�ы������BǄ�����x����,��� ǅ�����w��   9�0���t�������5  ��0���Q�f$ ���������������������������� ��������������������`�����������ƅ,��� ƅ%��� ������������������ ���������������������������0�����(����� ��������ǅ�����v������;�tU�8;�t@S�������� �G;�v	���sH�G�w����֍�����#��� ;�t
��j���ҋ�����P��  ���������  �������Q��4���Ǆ�����vPǅ4����v� ��������;�t*��h���Q������������RQP�JD  ������R��  ��������P��������������������  ��������;�t*��h���Q������������RQP��C  ������R�Y�  ��������P�������������������8�  �M���_^3͸   [�
 ��]� �������������U����  ��3ŉE��ESV��F �t��Q���   W�}j j	���Љ�t��Q���   j j���ЉF�t��Q���   j j���ЉF�t��Q���   j j
���ЉF�t��Q�J������P�у�������Rj������P���y-���t��Q�R�NQP�ҡt��H�A������R�Ћt��Q�J������P�ыt��B�P������Q�҃�������Pj������Q���-��P�������Bg  �������^$R���j  �������g  �t��H�A������R�Ћt��Q�J������P�у�h�r�������f  ������R���lj  �������Qg  �t��H�A������R�Ѓ�������Qj������R���c,��P�������f  �������~@P����i  ��������f  �t��Q�J������P�ыt��B�P������Q�҃�h�z��������e  ������P����i  �������f  j������V  ������Q���Jg  �t��R�Rhj h�   ������Q���ҡt��H�A������R�Ѓ�j@j������Q������?P  ��u+������J�������������y( u��j P��A  ��h��� �t��H�A�>  ������R�Ћt��Q�Jj j�������h�xP�ыt��B�P������Q�ҡt��H�Aj j�������hvR�Ѓ�(������Q������R���Gf  P������P������Q�C�����P������R�3���P� �t��H�A������R�Ћt��Q�J������P�ыt��B�P������Q�ҡt��H�A������R�Ћt��Q�J������P�у�$��l����8L  ǅl����v��l���R�� ��_^3�[�M�3��� ��]� ������R�Ћt��Q�Jj j�������h zP�ыt��B�P������Q�ҡt��H�Aj j�������h�zR�Ѓ�(������Q������R���	e  P������P������Q������P������R�����P�� �t��H�A������R�Ћt��Q�J������P�ыt��B�P������Q�ҡt��H�A������R�Ћt��Q�J������P�ы�����J��$j
������A  ��Ph�   ������Q�������T  ������:  ��u+������J�������������y( u��j P�	?  ������P�� ������>  �t��Q�J������P�ыt��B�Pj j�������hyQ�ҡt��H�A������R�Ћt��Q�Jj j�������hvP�ыt��B�P������Q�ҡt��H�Ij j�������R������P�у�<������R������P������Q������R�D�����P������P�4���P� �t��Q�J������P�ыt��B�P������Q�ҡt��H�A������R�Ћt��Q�J������P�ыt��B�P������Q�҃�$�~ ������P������������Q��������~ t-���   +��   ���Q���������t�������������������� j h  �� ����l�����H  ��l���Qǅl����v�A� �M���_^3͸   [�S ��]� ��������U��V��N+N��������������W�}�;�r�; �V����+�_��^]� �U��V��N+N���Q��������W�}�;�r��
 ��i��   F_^]� �����U��V��N+N��$I����������W�}�;�r�
 �V��    +�_��^]� ���������������U��V���U����Et	V�y�  ����^]� ��������������̡t�V��H�QV�����V ���   �V(R�V0�V8�V@�VH�VP�VX�V`�Vh�Vp�^x�t��H�A�Ћt��Q�J���   P�ыt��B�P���   Q�ҡt��H�A���   R�Ѓ���^át�V��H�A���   R�Ћt��Q�J���   P�ыt��B�P���   Q�ҡt��H�A���   R�Ћt��Q�BV�Ѓ�^��������U��V��V��v�� ���Et	V�?�  ����^]� �����U��A�U��Q �E��U+ЋA0�]� ��������������̋A �8 t�I0��3�����������������U��A�U��Q$�E��U+ЋA4�]� ���������������V���F@t�F�Q��  ���V�    �F �     �N0�    �V�    �F$�     �N4�    �f@��F<    ^������̍Q�Q �Q�Q$�A�A�Q(�Q0�A�A�Q,�Q4�     �A$�     �Q4�    �A�     �Q �    �A0�     ���������U��t�SV��H�QWV�ҡt��H�}�QVW���G�^���   �GS�^�G�F�O �N �W$�V$�G(�F(�O,�N,�W0�V0�G4�F4�O8�N8�W<�V<�G@�F@�OD�ND�WH�VH�GL�FL�OP�NP�WT�VT�GX�FX�O\�N\�W`�V`�Gd�Fd�Oh�Nh�Wl�Vl�Gp�Fp�Ot�Nt�Wx�Vx�G|�F|�t��Q�B�Ћt��QS���   P�J�ыt��B�H���   S�ыt��B�P���   SQ��ه�   ٞ�   �t��H�Q���   S�ҡt��H�A���   SR�Ћt��Q�B���   S�Ћt��Q�J���   SP�ы��   ��<_���   ��^[]� ��������U��VW�����u�E ���t��3ҋE����+��G����;Bw��t�	�3�;As� w��_^]� ���������U��VW�����u�� ���t��3ҋE�4�    +��G���;Bw��t�	�3�;As� w��_^]� ���������U��M����w3ɋ���+����R�n�  ����]Ã��3����xsڍEP�M��E    ��  h��M�Q�E�xv�J ���U��M����w3�i��   Q��  ����]Ã��3���=�   sߍEP�M��E    �  h��M�Q�E�xv�� ��������U��M����w3ɍ�    +���R��  ����]Ã��3����sڍEP�M��E    �=  h��M�Q�E�xv� ���U��EVP���i  �xv��^]� ����U��t�VW�}��H�QVW���G�^�G�^�G�F�O �N �W$�V$�G(�F(�O,�N,�W0�V0�G4�F4�O8�N8�W<�V<�G@�F@�OD�ND�WH�VH�GL�FL�OP�NP�WT�VT�GX�FX�O\�N\�W`�V`�Gd�Fd�Oh�Nh�Wl�Vl�Gp�Fp�Ot�Nt�Wx�Vx�G|�F|�t��Q�R���   P���   Q�ҡt��H�I���   R���   P��ه�   ٞ�   �t��B�@���   Q���   R�Ћt��Q�R���   P���   Q�ҋ��   ��(���   _��^]� ���U��S�]V�u;�t#W�}V���������   ���   ;�u��_^[]ËE^[]��������U��S�]V�u;�t#W�}���   ���   V���I���;�u��_^[]ËE^[]��������U��E��V��M�Q�F��v�P� ��V�H�N�P�V�@�F����^��]� ���������������U���E��QP� � ��]� ��������U��S�]V�u;�tW�y�WP��� �F��;�u�_��^[]� U���E��QP�� ��]� ��������U��S�]V�u;�tW�y�WP��� �F��;�u�_��^[]� U��E]� ������U��E�UV�1W��+�W�}WP�FR��_^]� �������������U��S�]VW�}��+�9us�= �E�MVSPQ�=� ����_^[]� �����������U��E]� ������U��E�UV�1W��+�W�}W�}WP�F(R��_^]� ���������U��S�]VW�}��+�9us�  �E�MVSPQ�� ����_^[]� �����������U��V��F��v��~�FP��  �}�NQ��  ���E��vt	V�R�  ����^]� �������̃��� ����������3��������������̃���������������U��U��@R�Uj�R��]� �������̋�� ������������ ������������̋A$�8 t�I4��3����������������̋A �8 t�Q0�: ~� � Ë�B�����V���P�҃��u�^ËF0��F ��Q��^����������U��E�p��3ɉH�H�H]� ���U��E�p��3ɉH�H�H]�  ���U��A � ��t<�Q;v5�U���t:P�t�A@u"�A0� �A ����t�A ����]� 3�]� ���]� ̋Q V�2��u���^�SW�y0����;�s�_[^��A@u/�A$� ��t&;�w9q<v9A<s�A<��A<+�I ��_[^�_[���^����������������U��SV�q$�W��t9A<s�A<�]����   �A �����   �E��u�A�y<+8�u��'��u��u�A�u��+8����t�5p���u����   �A� �y<+�;���   +Q0�)�Q ����   �Q$�����   �Q4�ЋA R��AR�R�����p��te���t_�E�=p���u�A�Y<+�u����u�A�u��+��	����u�u��|�A� �Y<+�;�+Q4�)�I$�
����5p��E_3ɉ0^�H�H�H[]� ��U��E�UVW�y$�4���t9A<s�A<�p�;���   S�]$��tR�Q ���tI��|w�A� �y<+�;�d+Q0�)�Q ��tX�Q$���tO�Q4�ЋA R��AR�R�����4��t-�?��t'��|#�A� �Q<+�;��Q4+��)�I$��p���[�E3�_�0�H�H�H^]�  ��������������U��V�q���Q�F�D��vP� �v��� ���Et	V���  ����^]� ����U��V��W�~8��v��t��襟��W���  ���N��� �Et	V��  ��_��^]� �������������U��V��W�w������~8��v��t���J���W�t�  ���N�}� �Et	V�]�  ��_��^]� ��U��Q�U�E�M���u	;A��   SVW�y;�st+�;�wn�   +���yr
���M�	����M��E�WQS�� ������t5�U�ERPV话������t,�M�+ލ|�WR�^S�a� ������u�_^���[��]� �E��x�Mr�	_��^+�[��]� �U��SV�uW��9ws�Q� �G+Ƌu;�s���]��;�r�Ãr�����MP�EP�W��������u;�s
_^���[]� 3�;���_^[]� �U��M����w3�Q��  ����]� ���3����s�EP�M��E    �� h��M�Q�E�xv��� �������������̋A �8 t�Q0�: ~����I ��P�� Ë�P���������V�����t(��u�� ��xr�H��H�@�9Fr�e� �F^����������U��E��u&�yr�I�E�U�]� �E�U���]� �yr�I����UP�EP�Q� � ��]� ���������U��QS��V�K��v��� j���  ������t@W�� ��A� j �M����Y� �G���s@�G�M��m� _�ˉs8�B���^��[��]�3��ˉs8�.���^��[��]�������U��S�]V�uW���    ��t)��t%�V�F��r����;�w��r� �N�;�v�1� �7�_��_^[]� ������������U��E�M�UV�uPQRV�� ����^]����������������U��E�M�U ��E��   ]� ����U��E�M��   ]� ������������U��E+E�M;�s��]� ����������U��S�]V�u��+θ����������������+ȋE�ȉM��;�t#+�W��I �<���x�   �;�u�E_^[]�^��[]����������������U��W�}��tV�u�   �^_]� ����U��M��t	�EP�����]� ���������U��S�]V�u��+˸����������������+���ɋыM��+�;�t+�W�M��M��x�<�   ���;�u�_^[]����������������U����US�]V�uW�}2��E��M��E��E�PQRWVS�r���+���Q���������i��   ����_^+�[��]����������U��j�h@fd�    PQSVW��3�P�E�d�    �e��E�    �]�}�u��$    ;utVW��������x�}��x�u���E������ǋM�d�    Y_^[��]�j j �� ����������������V��F � ��t=�N0�	��~�F0��F � �V �� ^Å�t�N0�9 ~����F ��Q���	��P���҃��u�^ËF �8 t�N0�9 ~��^Ë�P��^������U��QV3�9uW���u�~nS�]���������~6�M;ȋ�}��G ��UVQRS��� �G0)0u�)u�G ރ�0�u����P���҃��tF�C�M�u��} �[_��^��]� _��^��]� ������U��QV3�9uW���u�~mS�]���s�����~3�M;ȋ�}��VSP�G$�Q�<� �G4)0u�)u�G$ރ�0�u����P�B���Ѓ��tFC�M�u��} �[_��^��]� _��^��]� ������̋A��PV�q��D
��wW���w� ����~8��v��t���l���W��  ���N�� �F��H_�D1��v^�����������U���V���F@Wt �~$���t�N<;�s�F4� +��N4��E���u
_3�^��]� �V$�:S��t$�N4����;�s�	�v$�[�Q�_�^��]� �F@u=��u3���F4�N�+ߋ���� s�    ���v������+�;�s��u��u[_���^��]� �P�ND�E��������F��M���vSQ�M�QW�y����M�����u"�V�~<�:�F$�8�V4�E���F@u7�GPW�V�F$��+�V<� �V��+�+��V$ǉ��+�U��F4��F@t�V�:�F �     �V0�:��F$��F BR�+��RW��������M��F@t	Q���  ���F4�N@��v$��A��E[_�^��]� ������������U��S�]V��W9^s�� �F�}+�;�s����v^�N��r�V��V�U��r�V��V+�P�E��P+�Q�R�� �F+ǃ��~�Fr�N_� ��^[]� �N� _��^[]� ��U��} VW�}��t'�~r!�FS���vWSjP�� ��S���  ��[�~�F   �D> _^]� ����U��E�MPQ�� 3҃������]�V��~L t#��Pj��҃��t�FLP�t� ����}���^�3�^�U��A � S�]��t,�Q9s%���t�@�;�u�A0� �I �	��@���#�[]� �AL��t$���t�y< u��PQ�� �����t��[]� ���[]� �V��F ���t�Ћ�V0��;�s�^Ë�PW���ҋ����u_�^Ë�PW���ҋ�_^������������U��V��NLW��tl�U�}��u	��u�G�3�WPRQ��� ����uG�~L���FH�FA�<�����t�G�F�F�G�~ �~$�F0�F4�~L�`��FD_�F<    ��^]� _3�^]� ��������������U��ES�]V���F<    �F@����   ��<tzWS�ND��������ESPSW�� ���F@��F<u�N�9�V �:�N0��N@��u7��u�ǋV�:�N$���+ЋF4Ӊ�N �9 u�V�:�F �     �N0�9�N@_^[]� ����������U��V�1W�y��u�� 3��Mi��   �;xw��t�����3�;xs�Z� �E�x_�0^]� �����U��j�h`fd�    P��SVW��3�P�E�d�    �e����}�E�������v���"�_���鸫�������;�s�����+�;�w�4�E�    �NQ�������؉]��E������0�e��E�E�E�@P�M������E��E�   ��Ë}�u�]�M��v �r�G��GQP�VRS�� ���M�r�GP�W�  ���M�G�  ��w�O��r��� �M�d�    Y_^[��]� �u�~r�NQ��  ���F   �F    �F j j �� ����U����US�]V�uW�}2��E��M��E��E�PQRWVS�����+���Q���������i��   ���_^[��]��������������U��E�U;�tS�]VW����x�   ���;�u�_^[]�������U��V�uW�};�tS�]S����������   ;�u�[_^]�������U��j�h�fd�    PQSVW��3�P�E�d�    �e��E�    �]�}�u��$    ��v�EPV�������O�}��x�u���E������M�d�    Y_^[��]�j j ��� ��U��j�h�fd�    P��SVW��3�P�E�d�    �e��}�}��E�    �]�u��;utVW���r������   �}���   �u���E������ǋM�d�    Y_^[��]Ëu�};�t���R������   ;�u�j j �&� ���������������V��~r�FP���  ��3��F   �F�F^�����������U��VW�y��wP�������V��v�p� ���Et	W��  ����_^]� ��������U��yr�AV�uQP��������^]� V�u�AQP���������^]� ���������U��V���U����E3��w�u�   �u���t���t���E�x�Pr�@QRP���������^]� Q��RP��������^]� ��������U��U��V�p�d$ �@��u��M+�P�ARPj �'��������^]���������������U��Q�M�U�E� �E�P�EQ�MR�UPQR��������]�����U��Q�M�U�E� �E�P�EQ�MR�UPQR���������]�����U��j�h�fd�    P��SVW��3�P�E�d�    �e��u�u��E�    �]�}����v�EPV��� ���O�}���   �u���E������M�d�    Y_^[��]Ëu�};�t����������   ;�u�j j �� ���̃y$r�AÍA���U��V���,x�~$r�FP�u�  ��3��F$   �F �ΈF��� �Et	V�P�  ����^]� ������U��V���8x�~$r�FP�%�  ��3��F$   �F �ΈF�q� �Et	V� �  ����^]� ������U��SV3�S���� �^�   �F�^�F8�^4�^$�FT�^P�^@�Fp�EP�^lV�^\�� ����^[]� ���SV��WV�� ���~pr�F\P��  ��3ۿ   �~p�^l�^\�~Tr�N@Q�a�  ���~T�^P�^@�~8r�V$R�F�  ���~8�^4�^$�~r�FP�+�  ���~�^_�^��^[��� �����U��S�]V�����+F;�w�� ����   W�~����v�}� �F;�s9�NQW��������vZ�U�FRSP���h����~�~r:�F�8 _��^[]� ��uщ~��r�F_�  ��^[]� �F_�  ��^[]� �F�8 _��^[]� �����U��S�]VW�}��9_s�� ��E+�;�s���M;�uj��W���g���Sj ���]���_��^[]� ���v�� �M�F;�s�FPW�������M��vj�yr/�I�-��u�~��r�F_�  ��^[]� �F_�  ��^[]� ���~�^r���ËUW�Q�NQP�� ���~�~r��; _��^[]� ����������U��USVW���tF�~�F��r����;�r1��r���ȋ^�;�v��r� �MQ+�RV�������_^[]� �}���v�� �F;�s�VRW��������vY�N�^��r.��,��u�~��r�F_�  ��^[]� �F_�  ��^[]� �ËUWRQP��� ���~�~r��; _��^[]� �����U��Q�UV�uW�}�E� �E�P�ER��QPVW�9����΃���+΍�_^��]� ����U��V3���j��F�F   P�F�EP�������^]� ��������U���D��3ŉE��A �8 �M�t/�Ћ�Q0��;�s �A0��A ��Q���M�3��� ��]ËAL��u����M�3��� ��]Ãy< uP�� �����t����M�3��� ��]�SVWP�E�   �E�    �E� �U� ������  ��Pj�M��U����}��E���A  ���u؅�t!�ȃ�s�M�;�w�ȃ�s�M�U��;�v�.� �}��U�E�M����t�ȃ�s�M��;�r�� �}��U�E�ڃ���   ����t�ȃ�s�M�;�w�ȃ�s�M��;�v��� �}��U�E�M����t��s�E��;�r�� �}ЋO<��R�E�P�E�P�E�P�E�P�E��PV�GDP�҅��   ��~k����   �}���   j�U�R�M�����������P�E�jP�M� �u߃��M��(���_��^[�M�3���� ��]ÍM�M؋������u������E�9E���   �U��E����   ����t!�ȃ�s�M�;�w�ȃ�s�M�]��;�v��� �U��E�M����t��s�E�U��;�r�� �E�+�Pj �M�������OLQ�S� ������ ����M��h���_^���[�M�3��=� ��]Íu��m����}�M�Q�M�����������+}ԋ����~�UЋBL�M��T�NPR��� ������uߍM������M�_��^3�[��� ��]����������������U��V�u��W�x�I �@��u�+�PV�P���_^]� ����������U��SVW�}���    ��t�E9Fw;Fv�� �E�]���G9^w;^v�t� �]����t;�t�`� �O;�t!�F�E �UR�UR�URQPS�������F��_^[]� ��������U���,��3ŉE��y< �M���  �yA ��  ��Pj��҃��u2��M�3���� ��]ù   3��E� �M��E�E��E�   ��s�E�SV�@ W�E�U����  �؉]؅�t!�ȃ�s�M�;�w�ȃ�s�M�u��;�v�z� �U��E�M����t�ȃ�s�M�u��;�r�T� �U��E�}����   ����t$�ȃ�s�M�;�w�ȃ�s�M�]�ˋ]�;�v�� �U��E�M����t��s�E�U��;�r��� �E܋H<��R�E�P�E��SV��DP�҃� t<��t>���M��R  ����_^2�[�M�3��� ��]Í]�]�������u��V����E��@A �U��E����   ����t!�ȃ�s�M�;�w�ȃ�s�M�}��;�v�P� �U��E�M����t�ȃ�s�M�}��;�r�*� �U��E�}�+�tv����   ����t!�ȃ�s�M�;�w�ȃ�s�M�]��;�v��� �U��E�M����t��s�E�U��;�r��� �E܋HLQWjV�=� ��;�u7�U��E�M܀yA t0�������Wj�M��t���������u������u��h����M������M��_���_^�[�M�3��5� ��]ËM�3Ͱ�%� ��]�������������U��V�uW�};�t����I������   ;�u�_^]� ���������U��Q�UV�uW�}�E� �E�P�ER��QPVW������i��   ���_^��]� ����U��Q�U�E� �E�P�ER�U��Q�MPQR��������]� ��U��V�u�~r�FP�z�  ��3��F   �F�F^]� ���U��S�]V�u;�t!W�}j�j V�����������;�u��_^[]ËE^[]����������U�����3ŉE����M;�tT�PS�XV�p�]��YW�x�X�Y�X�Y�X�Y�X�Q�U��q�q�y�Q�P�p�q�Q�P_�p^�Q[�M�3��� ��]� ���U��V���9� 3��N�,xj��A�A   P�A�EP������^]� ����������U��V����� 3��N�,xj��A�A   P�A�EP������Dx��^]� ����V���,x�~$r�FP��  ��3��F$   �F �F��^�S� ��������������U��V�u3�j��NQ���F   �NP���Z�����^]� ���U���   SW�}3ۉ]���tm9uiVj荺  ������t)�Mj �E�P�   ����P��l����u���P��������3��^��t��l������������t�}�r�M�Q�/�  ��_�   [��]��U��V���� 3��N�8xj��A�A   P�A�EP�����Px��^]� ����V���8x�~$r�FP�Ȼ  ��3��F$   �F �F��^�� ��������������U��UV���W�F   �F    �F �x�@��u�+�PR�������_��^]� �����U���4��3ŉE�S�]�щU܃��u3�[�M�3��� ��]� �J$�9 Vt/�B4�	�0�;�s"��B$��Q��^��[�M�3���� ��]� �BL��t�z< u'P��P�� �����u�^���[�M�3��� ��]� �   3��E� �]؉M��E�E��E�   ��s�E��@ W�E�U������  �؉]ԅ�t!�ȃ�s�M�;�w�ȃ�s�M�u��;�v�_� �U��E�M����t�ȃ�s�M�u��;�r�9� �U��E�}����  ����t$�ȃ�s�M�;�w�ȃ�s�M�]�ˋ]�;�v��� �U��E�M����t��s�E�U��;�r��� �E܋H<��R�E�P�SV�E�P�E�P�E�P�E܃�DP�҅���  ���A  �U��E���"  ����t!�ȃ�s�M�;�w�ȃ�s�M�}��;�v�`� �U��E�M����t�ȃ�s�M�}��;�r�:� �U��E�}�+�tz����   ����t!�ȃ�s�M�;�w�ȃ�s�M�]��;�v��� �U��E�M����t��s�E�U��;�r��� �E܋HLQWjV�M� ��;���   �U��E�M��AA�M�9M���   �������}� �M���   j j�k���������]�]�������u��I����u�������u��<�����uu�U܋BL�M�PQ�^�������t �u�M��,���_��^[�M�3��� ��]� �M��������_��^[�M�3���� ��]� �M�������E_^[�M�3���� ��]� �M�������M�_^3̓��[�� ��]� �����������U���SV��F W�~@98u�}u�~< u�]K��]�~L ��   �W�����tw��u�}t�M�VLQSR�e� ����uX�NL�E�PQ�Y� ����uD�V 9:u�N�9�V �FA�Ή�V0+ȃ�A�
�E�M��U�_�H�ND^�     �P�H[��]� �E�p�_3�^��H�H�H[��]� �������������U����EV��~L �MW�}�E��M���   ��������t�FL�U�RP�$� ����uk��t�NLjWQ�� ����uT�FL�U�RP�|� ����u@�M�V �ND�N@9
u�FAPPQ�������E�M��U��H�ND_�     �P�H^��]�  �E�p�_��@    �@    �@    ^��]�  �����������U��QSVW�}���    ��t�E9Fw;Fv��� �E�]���G9^w;^v�� �]����t;�t�� �G;�tB�VPRS�����؋F���E���;�t��I ���������   ;}�u�E_�^^[��]� ��_^[��]� ����S��V�s3�;�t(W�{;�t���T������   ;�u�CP��  ��3�_^�C�C�C[����������������SV��3�W��9^Lt������u3��FLP�� ����t3��Έ^H�^A�h����^L�`���_�^<�ND^[����U��VW�}W���� 3�j��N�,x�GR�A   �QP�Q����_��^]� ����U���DSj3�hXx�M��E�   �]��]�������M���� j�S�E�P�M��E�,x�E�   �]܈]�����hH��M�Q�E�Dx�� �����������U��VW�}W����� 3�j��N�,x�GR�A   �QP�Q�\���_�Dx��^]� ��������������U���SVWj �M��5� �=4� �d��]�u+j �M��� �=4� u�0�@�0��4��M�� � �}�54��;ps"�H����u�x t诼 ;ps�P�4��3�����u]��t�M���ֻ _��^[��]ÍE�WP�C��������uhlx�M��f� h���M�Q��� �u��Ή5d��t��V�� ���M��� _��^[��]�������U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U���   SW�}3ۉ]���tp9ulVj�M�  ������t,�M�E�P�   �S���P��l����7����F    �Tw�3��7^��t��l�������`�����t�}�r�M�Q��  ��_�   [��]���������������U����US�]V�uW�}2��E��M��E��E�PQRWVS�B���+�$I�������������    +ȍ�_^[��]��������U��V�uW�};�t*S3ۃ~r�FP�O�  ���F   �^�^��;�u�[_^]����U��M3�;�tj��A�A   P�A�EP����]� �������U��j�h�fd�    P��SVW��3�P�E�d�    �e��}�}��E�    �]�u��;utVW���������}���u���E������ǋM�d�    Y_^[��]Ëu�};�t�]V���������;�u�j j �{� ����U��E���A�I��D#���   �} t	j j �N� ��t'h�x�M������E�P�M������h0��M�Q�"� ���M�t$h�x�Y����U�R�M������h0��E�P��� hxx�5����M�Q�M�����h0��U�R��� ��]� �����U��VW�}W���� 3�j��N�8x�GR�A   �QP�Q����_��^]� ����U��VW�}W���h� 3�j��N�8x�GR�A   �QP�Q�����_�Px��^]� ��������������U��QS3�V��WSS�^$�^�^�F  �F   �^�^�^ ����j��  ����;�t6�/� ��V� j �M����n� �C���s@�C�M�肷 �~$_^[��]�_�^$^[��]���������������U��V��~H ��wt����W�~8��v��t���4p��W�^�  ���N�g� �E_t	V�F�  ����^]� ������������U����A$SVW�8j �M��}�轶 �G���s@�G�M��Ѷ �M�Q�X�����j �M���葶 �G��v	���sH�G�w����֍M�#�薶 ��t
��j���Ћ�E�RP����_^[��]� ��U��V3�W�}��F�F�F;�u_2�^]� ��I�$	v����PW��������    +ύ��F�F_�V�^]� �����������U��j�h gd�    P��   ��3ŉE�SVWP�E�d�    �e��ًC��u3���K+ȸ���������������} �i  �s��p�����+K��������������º"""+ЋM;�s�L����;��,  ����"""+�;�s3���;�s��j W��������ȉ�p����u+s����������������E�    �EP�UR����+ƍ�Q������ǅl���   ��p���R�EP�KQ���Z���ǅl���   �U����+Ƌ�p�����R�CP�MQ���+����E������s�K+θ��������������E��t	V輫  ������+ϋ�p����ȉS�M����+эЉK�C�  ��p���R肫  ��j j �� ��+M��������������¹   �u��t����;E��   �}����+�����E�Q��p���RP���_����E�   �K��t���P+M���������������+�W�CP���Z����E�����s�[��t���R+�S�EP�:������N�E����+������p�����+�PPW��������C��p���QW�UR�������t���P�E�VP��������M�d�    Y_^[�M�3��D� ��]� ���������U��j�h0gd�    P���   SVW��3�P�E�d�    �e���u�F��u3���N+ȸ��Q��������ڋ}����  �N��+V���Q��������º�G+�;�s�h����8;��g  �����G+�;�s3���;�s��j S�j������ȉM�U+V���Q��������E�3҉U��U��URWi��   �P���[����E�   �E�P�MQ�VR�������E�   �E��i��   E�P�NQ�UR���|����E������N�V+Ѹ��Q������������t�VRQ�������FP��  ��i��   �E�؉^i��   ��~�F�M�d�    Y_^[��]� �]��u�}��~��i��   �QW�M��\�����~ �U�i��   �Pi��   �V�M��8���W�b�  ��j j �m� +M���Q���������;ύ������   �UR�;�����i��   �E�Q�VRP���p����E�   �N�����P+M���Q���������+�W�FP��������E�����^�v�����R+�V�EP�]������p�Ei��   �M�Q�R�U�P�k���j j �� �EP虽���^i��   ��+ǉESSP��������FS�MQ�UR����������P�E�WP�������������m����M�d�    Y_^[��]� ���������U��Q�M�U�E� �E�P�EQ�MR�UPQR�+�������]�����U���SVWj �M�腯 �=l� �h��]�u+j �M��i� �=l� u�0�@�0��l��M��p� �}�5l��;ps"�H����u�x t��� ;ps�P�4��3�����u]��t�M���&� _��^[��]ÍE�WP����������uhlx�M��� h���M�Q�7� �u��Ή5h��`g��V�S� ���M��Ϯ _��^[��]�������U��V�uW�};�tS�]j�j S���q�����;�u�[_^]������U��j�hPgd�    P��SVW��3�P�E�d�    �e��u�u��E�    �]�}����v�EPV���@���O�}���u���E������M�d�    Y_^[��]Ëu�};�t�]V��������;�u�j j �=� ������U��E�MP�����]����������������U��U��t�Ay( u���URP�~���]� ���������̋A��PV�q��D
��x�~H W��wt�������~8��v��t���ff��W萤  ���N虱 �F��H_�D1��v^�����U��EVWP���p�������B�����Є�t�G<    _^]� �ωw<����_^]� �U���   ��3ŉE�SV�ًCW�   �u�}��{�u��+ȸ��������������;�vH9{v��� �K+K�E�P���������������+�VWP���r���_^[�M�3�芸 ��]�| s]9{v�� �K���t����M�;Kv�� �M���M�V��|�����|���������t����M���|���WPQR��t���P�������M�_^3�[�� ��]�| �������������U���SV��^�F��+ȸ��Q��������W�}�;�vD9^v��� �V+V��EP���Q���������+�WSQ���p����M����_^[��]�� sN9^v�� �F��M��E;Fv�� �E��E�W�E�P�M��U�������M��P� SQRP�M�Q���o����M臶��_^[��]�� ��������������U��E�UP��Q�MQR������]� �U��V��~L W��   �E�M�UPQR�� ��������   ���FH�FA 蒷���N8�G�F�F�G�~ �~$�F0�F4�~L�`��FD�F<    �9j �M�}�N� �G���s@�G�M�b� �UR��������P�����҄�t�M�F<    �8c��_��^]� �Ή~<�����M�c��_��^]� _3�^]� ��������������U��Q�U�E� �E�P�ER�U��Q�MPQR��������]� ��U��j�hpgd�    P��0��3ŉE�SVWP�E�d�    �e��}�u�ủu��E�   3��E�EԉE��]�;}t$�E�PV���o���WV�x��������ũ��}����E������}�r�M�Q�q�  ���ƋM�d�    Y_^[�M�3��9� ��]Ëuȋ}�;�t�]�I V��������;�u�3�PP�?� ��������V���HW�13��@u�@(��ȋB0�Ѓ��u�   ��I΅�t�Aǃy( u��j P�u���_��^�U��QV��F��t�M�Q�N�VRQP�@����VR觟  ���P�F    �F    �F    臟  ��^��]����������������U��VW�y��wX������V��v�� ���Et	W�C�  ����_^]� ��������U��j�h�gd�    P��SVW��3�P�E�d�    �e���u��H΋A����   �I,��t������} up��P�L2��tb�MQ����1a��P���������M�~`���E�    ��B�L0(�����E���uj j��I�������ЋG�PHu+�E�������Q�2�y ue��M�d�    Y_^[��]� ��Q�L2(�����럋M��@��H���x( u�����H�Hu�E������I9Ëu��j j �� �A���y( u��j P����2��M�d�    Y_^[��]� ������������U��SVW�}���    ��t�E9Fw;Fv蠻 �E�]���G9^w;^v脻 �]����t;�t�p� �O;�t5�F�E �UR�UR�URQPS�w����V�؋EP�NQRS�������(�^��_^[]� ����U��Q�UV�uW�}�E� �E�P�ER��QPVW�9�������    +΍�_^��]� ��U��SV�uW�}��+ϸ�$I�����������    +ȋE�ɋ�+�;�t+ƉE��E��V�0�o���;�u�_^��[]�����U���SV��FW�E�9Fv�l� �~�;~v�]� �M��QSWP�U�R������_^[��]������������U��QS3�VW�ىE�9Et��x�CX�v��Q��v�C��p��������{j �Ή~(�F,    �����~( �F0u�F��j P���d����F    ��Q����x��������w�GH �GA �E���3��GL�`��G<�OD_^��[��]� ���������U��QS3�VW���E�9Et��x�GP�v��Q��v�G��p��������_j �Ή^(�F,    ������~( �F0u�F��j P�������E�F    ��Q�M��PQ����w������_^[��]� ����U��j�h�gd�    P��SVW��3�P�E�d�    �e���u�3ۉ]�^�u܋�H�D1(;�t�H諧 j���G�����tY�}��~R�E�    ��B�L0(觸���E���u���&�M;�u�F��Q�L2(�q����O�}��m���]��E������E�  �~ u���Ӌ�I΅�t�Ay( u��j P�����E܋�J�D(��t�H�� �ƋM�d�    Y_^[��]� �F�M�A�M��H�L1(�0����D����M��B��H���x( u�����H�Hu�E�������=Ëu�]��E���j j �m� ������U��j�h�gd�    P��$SVW��3�P�E�d�    �e�3��}��E� �u�uЋ�H�D1(��t�H�,� j �����������   ��BƋ@$�8�}�j �M��� �G���s@�G�M�蓡 �E�P�������E܍M��|Z��j�j �]��������E�    ��Q�2�A��~���r��������}؋I(������E��v	���uq�M��E������}��H�D1    �}� u����J΅�t�Aǃy( u��j P������EЋ�Q�D(��t�H�<� �ƋM�d�    Y_^[��]��ȋU܋R�JHu�Pj��������E�O�}؋�H�L1(�U����O����M��B��H���x( u�����H�Hu�E�������?Ëu�-���j j 蕵 ��������������U��Q�U�E� �E�P�ER�U��Q�MPQR�K�������]� ��U��Q�M�U�E� �E�P�EQ�MR�UPQR�;�������]�����U��QVW�}��;��W  �G�O+ȸ�$I����������Eu���V���_��^��]� �NS�^+˸�$I�����������9MwY�GSP�GP�}����MQ�N�VRQP�����O+O��$I�������������    +ЋF[��_�N��^��]� ��u3���V+ӉU���$I���U��������9Ew+�G��    +э�SQP�M������F�O�U��PQR�M��t�FPS�������FP��  ���O+O��$I�����������P���!�����t�N�W�GQRP���z����F[_��^��]� ������������U��j�h hd�    P��<��3ŉE�SVWP�E�d�    �e���u��E�E��F��u�E���N+ȸ�$I����������E̋}����  �^��+N��$I����������¹I�$	+�;�s����ǋM�;���  ����I�$	+�;�s�E�    �M��ʉM�;�s�E̋�j Q�������ȉMȋ]+^��$I����������ډ]�3��E��E��U�RW��    +Í�Q���W����E�   �U�R�EP�NQ��������E�   ߍ�    +ӋEȍ�Q�VR�EP��������E������^�N+˸�$I��������������t�VRS��������FP���  ���E̍�    +ȋEȍ��V��    +ύ��V�F�  �]��uċ}ȃ�~��    +ƍ�QW�M��e�����~(�U���    +ȍ�R��    +ƍ�Q�M��9���W�s�  ��j j �~� +]��$I�����������;���   �M�Q�M��������    +��ۋE�R�NQP�������E�   �N�U�R+M��$I�����������+�W�FP��������E�����^�v�M�Q+�V�UR��������~�M��    +����M��Q�R�U�P�e���j j 賰 �E�P�M��@����F�Eč�    +��ۋ�+�PPW��������F�M�QW�UR�����E�P�E�SP�^������M��C����M�d�    Y_^[�M�3��� ��]� �����U��EV���F�@   �@    �@ ���t#PQ������Q���D��t�    ^]� ��^]� U���SV��^W�~��+ϸ�$I�����������u3��3;�v蠯 �M���t;�t莯 �M+ϸ�$I������������M�U�EQjRP��������^;^v�T� �6W�M��u��]��L����E�M��U�_^��P[��]� �����U���SVW���G��u3���O+ȸ�$I�����������_��+O��$I�����������;�s.�U�E� �M�Q�MR�GPQjS����������__^[��]� 9_v袮 �U�RSP�E�P������_^[��]� ���������������U��EW�};E,tQ���u�^� �ML�EP�+����E��u�F� �E��t#�MQP�������J���Dt3��E��E;E,u��}(�UL�r�EP���  ���}H�E(   �E$    �E r�M4Q�؏  ����_]�U��QSV�u3ۈ]��E��M��U�P�ELQ�M,RP�� �ĉj��HS�U0�A   �YR�Y�,����M�� �ĉj��HS�U�A   �YR�Y����V�������T�}(r�EP�N�  ���}H�E(   �]$�]r�M4Q�/�  ����^[��]�����U��p���t]��]���������������̡t����   �p�ǀ�   0H�p   �������������������������������U��E�� t��t3�]ù���7 �����]ø   ]����j j j jdjdhZ� j���w*  � ����U���VWh{jh��jH��  ������t���u< �N��z������3��t��H�A�U�R�Ћt��Q�Jj j��E�h {P�у��U�R�M��hB �8Vj��, ��PWj j��, ��PhZ� �> ���M����UC �t��H�A�U�R�Ѓ�_��^��]����������U��V��N�R�������; �Et	V��  ����^]� ��%p�%p�%p�%p������������U��E�t�� ]��U��t��P�EP�EP�EPQ�J�у�]� �����������̡t�V��H�QV�ҡt��H$�QDV�҃���^�����������U��t�V��H�QV�ҡt��H$�QDV�ҡt��U�H$�AdRV�Ѓ���^]� ��U��t�V��H�QV�ҡt��H$�QDV�ҡt��U�H$�ARV�Ѓ���^]� ��U��t�V��H�QV�ҡt��H$�QDV�ҡt��H$�U�ALVR�Ѓ���^]� �̡t�V��H$�QHV�ҡt��H�QV�҃�^�������������U��t��P$�EPQ�JL�у�]� ����U��t��P$�R]�����������������U��t��P$�Rl]����������������̡t��P$�Bp����̡t��P$�BQ�Ѓ����������������U��t��P$��VWQ�J�E�P�ыt��u���B�HV�ыt��B�HVW�ыt��B�P�M�Q�҃�_��^��]� ���U��t��P$�EPQ�J�у�]� ����U��t��P$��VWQ�J �E�P�ыt��u���B�HV�ыt��B$�HDV�ыt��B$�HLVW�ыt��B$�PH�M�Q�ҡt��H�A�U�R�Ѓ� _��^��]� ���U��t��P$��VWQ�J$�E�P�ыt��u���B�HV�ыt��B$�HDV�ыt��B$�HLVW�ыt��B$�PH�M�Q�ҡt��H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e����t��Q$�JH�E�P�ыt��B�P�M�Q�҃���^��]� ����̡t��P$�B(Q��Yát��P$�BhQ��Y�U��t��P$�EPQ�J,�у�]� ����U��t��P$�EPQ�J0�у�]� ����U��t��P$�EPQ�J4�у�]� ����U��t��P$�EPQ�J8�у�]� ����U��t��UV��H$�ALVR�Ѓ���^]� ��������������U��t��H�QV�uV�ҡt��H$�QDV�ҡt��H$�U�ALVR�Ћt��E�Q$�J@PV�у���^]�U��t��UV��H$�A@RV�Ѓ���^]� ��������������U��t��P$�EPQ�J<�у�]� ����U��t��P$�EPQ�J<�у����@]� ���������������U��t��P$�EP�EPQ�JP�у�]� U��t��P$�EPQ�JT�у�]� ���̡t��H$�QX�����U��t��H$�A\]�����������������U��t��P$�EP�EP�EPQ�J`�у�]� �����������̡t��H(�������U��t��H(�AV�u�R�Ѓ��    ^]��������������U��t��P(�R]����������������̡t��P(�B�����U��t��P(�R]�����������������U��t��P(�R]�����������������U��t��P(�R ]�����������������U��t��P(�E�RjP�EP��]� ��U��t��P(�E�R$P�EP�EP��]� �t��P(�B(����̡t��P(�B,����̡t��P(�B0�����U��t��P(�R4]�����������������U��t��P(�RX]�����������������U��t��P(�R\]�����������������U��t��P(�R`]�����������������U��t��P(�Rd]�����������������U��t��P(�Rh]�����������������U��t��P(�Rl]�����������������U��t��P(�Rx]�����������������U��t��P(���   ]��������������U��t��P(�Rt]�����������������U��t��P(�Rp]�����������������U��t��P(�BpVW�}W���Ѕ�t:�t��Q(�Rp�GP���҅�t"�t��P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U��t��P(�BtVW�}W���Ѕ�t:�t��Q(�Rt�GP���҅�t"�t��P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U��VW�}W���0�����t8�GP���!�����t)�OQ��������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W���0�����t8�GP���!�����t)�O0Q��������t��HW��������t_�   ^]� _3�^]� ������������U����t��E�    �E�    �P(�RhV�E�P���҅���   �E���uG�t��H�A�U�R�Ћt��Q�E�RP�M�Q�ҡt��H�A�U�R�Ѓ��   ^��]� �t��Qhx{he  P���   �Ћt����E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�  ��3�^��]� �M��U�j IQ�MR������E�P��~  ���   ^��]� ���������������U��t���V��H�A�U�R�Ѓ��M�Q������^��u�t��B�P�M�Q�҃�3���]� �t��H$�E�I�U�RP�ыt��B�P�M�Q�҃��   ��]� �U��Q�t��P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U��t��P(�R8]�����������������U��t��P(�R<]�����������������U��t��P(�R@]�����������������U��t��P(�RD]�����������������U��t��P(�RH]�����������������U��t��P(�E�R|P�EP��]� ����U��t��P(�RL]�����������������U��t��E�P(�BT���$��]� ���U��t��E�P(�BPQ�$��]� ����̡t��H(�Q�����U��t��H(�AV�u�R�Ѓ��    ^]��������������U��t��P(���   ]��������������U��t��H(�A]����������������̡t��H,�Q,����̡t��P,�B4�����U��t��H,�A0V�u�R�Ѓ��    ^]�������������̡t��P,�B8�����U��t��P,�R<��VW�E�P�ҋu���t��H�QV�ҡt��H$�QDV�ҡt��H$�QLVW�ҡt��H$�AH�U�R�Ћt��Q�J�E�P�у�_��^��]� �������U��t��P,�E�R@��VWP�E�P�ҋu���t��H�QV�ҡt��H�QVW�ҡt��H�A�U�R�Ѓ�_��^��]� ��̡t��H,�j j �҃��������������U��t��P,�EP�EPQ�J�у�]� U��t��H,�AV�u�R�Ѓ��    ^]�������������̡t��P,�B����̡t��P,�B����̡t��P,�B����̡t��P,�B ����̡t��P,�B$����̡t��P,�B(�����U��t��P,�R]�����������������U��t��P,�R��VW�E�P�ҋu���t��H�QV�ҡt��H$�QDV�ҡt��H$�QLVW�ҡt��H$�AH�U�R�Ћt��Q�J�E�P�у�_��^��]� �������U��t��H��D  ]��������������U��t��H��H  ]��������������U��t��H��L  ]��������������U��t��H�I]�����������������U��t��H�A]�����������������U��t��H�I]�����������������U��t��H�A]�����������������U��t��H�I]�����������������U��t��H���  ]��������������U��t��H�A]�����������������U���V�u�E�P��������t��Q$�J�E�P�у���u-�t��B$�PH�M�Q�ҡt��H�A�U�R�Ѓ�3�^��]Ët��Q�J�E�jP�у���u=�U�R��������u-�t��H$�AH�U�R�Ћt��Q�J�E�P�у�3�^��]Ët��B�HjV�у���u�t��B�HV�у����I����t��Q$�JH�E�P�ыt��B�P�M�Q�҃��   ^��]�����������U��t��H�A ]�����������������U��t��H�I(]�����������������U��t��H��  ]��������������U��t��H��   ]��������������U��t��H��  ]��������������U��t��H��  ]��������������U��t��H�A$��V�U�WR�Ћt��Q�u���BV�Ћt��Q$�BDV�Ћt��Q$�BLVW�Ћt��Q$�JH�E�P�ыt��B�P�M�Q�҃�_��^��]������U��t��H���  ��V�U�WR�Ћt��Q�u���BV�Ћt��Q$�BDV�Ћt��Q$�BLVW�Ћt��Q$�JH�E�P�ыt��B�P�M�Q�҃�_��^��]���U��t��H���  ]��������������U���<���SVW�E�    ��t�E�P�   �������/�t��Q�J�E�P�   �ыt��B$�PD�M�Q�҃��}�t��H�u�QV�ҡt��H$�QDV�ҡt��H$�QLVW�҃���t)�t��H$�AH�U�R����Ћt��Q�J�E�P�у���t&�t��B$�PH�M�Q�ҡt��H�A�U�R�Ѓ�_��^[��]���U��t��H�U���  ��VWR�E�P�ыt��u���B�HV�ыt��B$�HDV�ыt��B$�HLVW�ыt��B$�PH�M�Q�ҡt��H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]����������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]�������������̡t��H���   ��U��t��H���   V�uV�҃��    ^]�������������U��t��P�]��t��P�B����̡t��P���   ��U��t��P�R`]�����������������U��t��P�Rd]�����������������U��t��P�Rh]�����������������U��t��P�Rl]�����������������U��t��P�Rp]�����������������U��t��P�Rt]�����������������U��t��P���   ]��������������U��t��P��  ]��������������U��t��P�Rx]�����������������U��t��P���   ]��������������U��t��P�R|]�����������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P�EPQ��  �у�]� �U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��E��t �t��R P�B$Q�Ѓ���t	�   ]� 3�]� U��t��P �E�RLQ�MPQ�҃�]� U��E��u]� �t��R P�B(Q�Ѓ��   ]� ������U��t��P�R]�����������������U��t��P�R]�����������������U��t��P�R]�����������������U��t��P�R]�����������������U��t��P�R]�����������������U��t��P�R]�����������������U��t��P�E�R\P�EP��]� ����U��t��P�E��  P�EP��]� �U��t��E�P�B ���$��]� ���U��t��E�P�B$Q�$��]� �����U��t��E�P�B(���$��]� ���U��t��P�R,]�����������������U��t��P�R0]�����������������U��t��P�R4]�����������������U��t��P�R8]�����������������U��t��P�R<]�����������������U��t��P�R@]�����������������U��t��P�RD]�����������������U��t��P�RH]�����������������U��t��P�RL]�����������������U��t��P�RP]�����������������U��t��P���   ]��������������U��t��P�RT]�����������������U��t��P�EPQ��  �у�]� �U��t��P���   ]��������������U��t��P���   ]��������������U��t��P�RX]����������������̡t��P���   ��U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]��������������U��t��P���   ]�������������̡t��P���   ��U��t��P���   ]�������������̡t��P���   ��t��P���   ��t��P���   ��U��t��H���   ]��������������U��t��H��   ]��������������U��t��H�U�E��VWRP���  �U�R�Ћt��Q�u���BV�Ћt��Q�BVW�Ћt��Q�J�E�P�у�_��^��]������������U��t��H���  ]��������������U��t��P(�BPVW�}�Q�]���E�$�Ѕ�tM�t��G�Q(�]�E�BPQ���$�Ѕ�t,�t��G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U��t��P(�BTVW�}����$���Ѕ�tE�t��G�Q(�BT�����$�Ѕ�t(�t��G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U��t��P(�} �R8����P��]� �U��t��P�BdS�]VW��j ���Ћt��Q�����   hx{Fh�  V�Ћt����E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћt��Q(�BHV���Ѕ�t �t��Q(�E�R VP���҅�t�   �3��EP�g  ��_��^[]� ������U���V�E���MP�k���P���#����t��Q�J���E�P�у���^��]� ��̡t��P�BVj j����Ћ�^���������U��t��P�E�RVj P���ҋ�^]� U��t��P�E�RVPj����ҋ�^]� �t��P�B�����U��t��P���   Vj ��Mj V�Ћ�^]� �����������U��t��P�EPQ�J�у�]� ����U��t��P�EPQ�J�у����@]� ���������������U��t��P�E�RtP�ҋt����   P�BX�Ѓ�]� ���U��t��P�E�Rlh#  P�EP��]� ���������������U��t��P�E�RlhF  P�EP��]� ���������������U��t��P�E�RtP�ҋt����   �M�R`QP�҃�]� ���������������U��t��P���   ]��������������U��t��P�E���   P�҅�u]� �t����   P�B�Ѓ�]� ��������U���V�u�W�}�����Dz�F�_����D{:�F����$��� �G��$�]��� �E���������D{_�   ^��]�_3�^��]���������U���VW�M��`����E�}��t-�t��Q4P�B�Ѓ��M��u����_3�^��]Ë�R(��t��H0�QW�҃��M��tԋ�R Q�MQ���ҋ�t��P�B �M��Ѓ��t�t��Q0�Jx�E�PW�у��M��.���_��^��]�������U��t��P�B VW�}�����=NIVb��   ��   =TCAbtR=$'  t6=MicM��   �t��Q���   j hIicM���ЋWP�B����_^]� ��BW����_�   ^]� �t��Q���   j hdiem���ЋWP�B����_^]� =INIb��   �~ u���B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� �a�  _3�^]� =cnys����_3�^]� ������V����{�t��H0�Vh@o�҉F���F    ��^�����V��F��{��t�t��Q0P�B�Ѓ��F    ^�����̡t��P0�A���   P�у����������U��t��P0�E�I���   PQ�҃�]� �������������̡t��I�P0���   Q�Ѓ���������̡t��P0�A���   j j j j j j j j j4P�у�(������̡t��P0�A���   j j j j j j j j j;P�у�(�������U��t��P0�E�IPQ���   �у�]� ��������������U����E V��P�M��;����t��E�Q�R4Ph8kds�M��ҡt��E     �H0���   �U R�U�E�P�Ej R�UP�ER�UP�FRj2P�ыu ��(�M��������^��]� ��������������̡t��I�P0���   Q�Ѓ����������U��V��F��u^]� �t��Q0�M ���   j j j j j Q�Mj QjP�ҡt��H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uËt��Q0P�B�Ѓ������̋A��u� �t��Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5t��v0Q�MQP���   R�U�R�Ћu�    �F    �t����   j P�BV�Ћt����   �
�E�P�у�$��^��]� �������U��t��P0�E�I�RPQ�҃�]� �U��A��t)�t��Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5t��v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5t��v0QP���   R�Ѓ�^]� �����������U��Q��u3�]� �E�H� V�5t��v0Q�MQPR�V\�҃�^]� ����������U��A��u]� �t��Q4�M��  Q�MQP�҃�]� �U��A��u]� �t��Q4�M�RhQ�MQP�҃�]� ����U��A��u]� �t��Q4�M�RpQ�MQP�҃�]� ����U��A��u]� �t��Q4�M��  Q�MQP�҃�]� �U���$VW��htniv�M��I����t��P�E�R4Phulav�M��ҡt��P�B4hgnlfhtmrf�M��Ћt��E�Q�R4Phinim�M��ҡt��P�E�R4Phixam�M��ҡt��P�E�R4Phpets�M��ҡt��P�E�R4Phsirt�M��ҋE �}$=  �u�����t.�t��QP�B4h2nim�M��Ћt��Q�B4Wh2xam�M��ЋU�M�QR�E�P�������t����   P�B8�Ћt����   �
���E�P�у��M��h���_��^��]�  ��������������U���$V��htlfv�M�������E�t��P�B,���$hulav�M��Ћt��E,�Q�R4Phtmrf�M����E�t��P�B,���$hinim�M����E�t��Q�B,���$hixam�M����E$�t��Q�B,���$hpets�M��Ћt��ED�Q�R4Phsirt�M��������E0��������Dzw���]8����Dzm�؋t��E@�Q�R4Phdauq�M��ҋM�E�PQ�U�R���/����t����   P�B8�Ћt����   �
���E�P�у��M�������^��]�@ �١t��P�B,���$h2nim�M����E8�t��Q�B,���$h2xam�M����V�����U���$V��hgnrs�M��j����E�t��E��E�   �Q���   �E�Pj�M��ҡt����   ��U�R�ЋM�t��M����E�   �B���   �M�Qj�M��ҡt����   ��U�R�ЋU���M�QR�E�P�������t����   P�B8�Ћt����   �
���E�P�у��M��������^��]� �U���$V��hmnrs�M������t��P�E�R4Pj�M��ҋM�E�PQ�U�R�������t����   P�B8�Ћt����   �
���E�P�у��M��n�����^��]� �����U��E��$�����VDSSS��P�M�������t��Q�B �M��Ћt��QjP�B4�M��ЋU�M�QR�E�P��������t����   P�B8�Ћt����   �
���E�P�у��M��������^��]� �����������U���$V��hCITb�M��j����t��P�E�R8PhCITb�M��ҡt��P�E�R4Phsirt�M��ҡt��P�E�R4Phulav�M��ҋM�E�PQ�U�R���<����t����   P�B8�Ћt����   �
���E�P�у��M�������^��]� U��E��Vj ��P�M�Q�M������UPR���)�����t��H�A�U�R�Ѓ���^��]� ����������U��E,��UPj ���T$�$htemf�E$�� �\$�E�\$�E�\$�E�$R�/���]�( �����������U��� |�E��������{��{��D{����������{�E��������D{����E,��Pj ���T$�U�$hrgdf�E$�� �������\$���\$�\$�E�$R����]�( ���������U��E,��Pj ���T$�U�$htcpf�E$�� ��v�����\$�E���\$�}�\$�E�$R�C���]�( ���������������U��Q��u3�]� �E�E�H� V�5t��v0Q�M Q�M���\$�E�$QPR�V(�҃�$^]� ������U��Q��u3�]� �E�H� V�5t��v0Q�MQPR�V,�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5t��v0Q�MQPR�V,�҃�^]� ����������U��Q��u3�]� �E�H� V�5t��v0Q�MQPR�V0�҃�^]� ����������U��SVW���W��t$�E�H�5t��^0� �uQVP�C0R�Ѓ���u	_^3�[]� �W��t��E�H� �t��[0Q�NQPR�S0�҃���t̋W��tŋE�H� �=t��0Q��VP�G0R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5t��v0Q�MQ�MQPR�V<�҃�^]� ������U��QV3�W��u3��,�E�H� �5t��v0Q�MQPR�V,��3Ƀ�9M������t��M�B�P0VQ�M�ҋ�_^]� ����U��AV��u3��"�M�Q�	�5t��v0R�URQP�F,�Ѓ����t��Q�E�M�R4PQ�M�ҋ�^]� ���������������U��A��V��u3��"�M�Q�	�5t��v0R�U�RQP�F0�Ѓ����t��E��Q�E�M�R,���$P�ҋ�^��]� �����U�����V���U�V�U��]�W��t$�E�H� �=t��0Q�M�QPR�W0�҃���u
_3�^��]� �V��t�E�H� �=t��0Q�M�QPR�W0�҃���tˋV��tċE�H� �5t��v0Q�M�QPR�V0�҃���t��t��P�M�RH�E�PQ�M��_�   ^��]� �����������U��� ��A�U�V�U�W�]���u3��&�M�Q�	�5t��v0R�U�R�U�RQP�F<�Ѓ����E�}���t�t��Q�RH�M�QP���ҋE���t�t��E��Q���$P�B,����_��^��]� U��t��P�E���   Vj ��MP�ҋM$�U Q�MR�Uj Q�MR�UQPR������^]�  ����������U��t���P�E���   V���$��MP���E8�E@�M,�Uj P���\$�E0�$Q�E$�� �\$���E�\$�E�\$�$R�����^]�< ������U��t���P�E���   V���$��MP����Ej j ���T$���$htemf�E$�� �\$�E�\$�E�\$�$P����^]�$ �����������U��t���P�E���   V���$��MP���E$�Ej �� �\$���E�\$�E�\$�$P����^]�$ ��������������U��t���P�E���   V���$��MP����j j ���T$�E�$htcpf�E$�� ��v�������\$�E���\$�}�\$�$P����^]�$ ���������������U��t��� V��H�A�U�R�ЋM�E��Qj �U�RP�M�Q�M�����UPR���������t��H�A�U�R�Ћt��Q�J�E�P�у���^��]� ������������U���dV��M������t��Q���   P�EP�M�Q�M��P�M������M��Q���j j �E�P�M������MPQ���U����t����B�P�M�Q�҃��M������M�������^��]� �����U���P��EV�]���W�}����t�t��Q���$P���   �����]���t��U��UЍE��]؋Q�M���   PQ�E�P���ҋ�M��P�U�H�M�P�U�H�M��P�F�U��u_^��]� �M�E�Q�	�5t��v0R�U R���\$�U��E��$RQP�F(�Ѓ�$_^��]� ���������������U���0�E�M���u�t��H���   �҅�u��]� SVW���_  ��htlfv�MЉu�z����E�}�t��X�U�����$茂 �]��G�$�~� �}�S,�M��$hulav�ҡt��P�B4hmrffhtmrf�M��Ћ}��t��M�Y���$�5� �]��G�$�'� �}�S,�M��$hinim�ҋ}��t��M�X���$��� �]��G�$�� �}�S,�M��$hixam����t��P�B,���$hpets�M��Ћt��Q�B4j hdauq�M��Ћt��Q�B4Vhspff�M��Ћt��E �Q�R4Phsirt�M��ҋM�E�PQ�M��U�R�^����t����   P�B8�Ћt����   �
���E�P�у��M��;���_��^[��]� U��E��V���u�t��H���   �҅�u^��]� ���N]  �E�F��u3��"�M�Q�	�5t��v0R�U�RQP�F0�Ѓ����E���|�M������\$�M��$��	 ��M��P�Q�P�Q�@�A��^��]� ����������U���0��t��]�V���M�]�P���   �E�PQ�M�E�P�ҋ�P�M��Hj �U�P�E P�M��MQ�M�U��UR�U�E�PQR������^��]� ���������������U�����UV�]���E�P�]��ERP�����t��Q�M�R@���E�PQ�M�ҋ�^��]� ����������U��A��u]� �M�Q�	V�5t��v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� �t��Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� �t��Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U��t��P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� �t��Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj>P�ҋE���(��]� ������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5t��v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M��X �MQ�U�R�M�� ��tm�}��E��tN�t����   P�BH�ЋM��I����tQ�W�7�t��[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M��; ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5t��v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� �t��E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �t��Q0�M�RDQ�MQ�MQP�҃�]� U��A��u]� �t��Q0�M�RHQ�MQ�MQ�MQ�MQ�MQP�҃�]� ���̋A��uËt��Q0P�BX�Ѓ�������U��A��u]� �t��Q0�M�RLQ�MQP�҃�]� ����U��A��u]� �t��Q0�M�RP��   �QP�҃�]� ��U��A��u]� �t��Q0�M�RPQP�҃�]� ��������U��A��u]� �t��Q0�M�RTQ�MQ�MQ�MQP�҃�]� ������������U��t�V�u�VW���H4�R�ЋE�F    �~�H� �t��R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� �t��Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I�t��R0P�EPQ���   �у�]� ������̡t��I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u���� �t��R0�I�R@V�uVP�EPQ�҃�^]� �����������U��t��P0�E�I�RdP�EP�EP�EP�EPQ�҃�]� �U��t��P0�E�I�RpP�EP�EP�EP�EPQ�҃�]� �U��E�P� V�5t��v0R�UR�UR�UR�URP�A�NhP�у�^]� ��������U��E� �t��R0j j j j j j j P�A���   jP�у�(]� �����������U��E� �t��R0j j j j j jj P�A���   jP�у�(]� �����������U��E� �t��R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M������E�H� �t��R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R������M�������^��]� ����������U��E�P� V�5t��v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5t��v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5t��v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5t��v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U��t��P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U��t��UVj j j j j R��H0�E�Vj P���   jR�Ћt��Q0�E�N�RtPQ�҃�0^]� ��U��t��P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡t��P0�A���   j j j j j j j j jP�у�(�������U��t��P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡t��P0�A���   j j j j j j j j j(P�у�(�������U��t��P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U��t��P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡t��P0�A���   j j j j j j j j jP�у�(������̡t��P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}�M���t�t��P���   j j���Љ�u��t�t��Q���   j j���Љ�t��Q0�E��H�R`VWQ�҃�_^[��]� �U��t��P0�E�I���   P�EP�EPQ�҃�]� �����̡t��P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V����{�t��H0�Vh@o�҉F3��F�F���|�F   ��^�������V��F��{��t�t��Q0P�B�Ѓ��F    ^������U��E�UVj ��MP�EQ3�9MR��Pj �F    ��
Q��������t�~ t
�   ^]� 3�^]� �U��E�A�I��u3�]� �t��B0Q�H�у�]� ����U��t��P�B S�]V�����=ckhc��   ��   =cksate=TCAb��   �t��Q���   Wj hdiem���Ћ���BSW���F   �Ѓ~ ��t��t��u3Ƀ���Q���C���_^��[]� �~ tK��B����^[]� �~ t6��������t+�F    ^�   []� =atnit�MQS������^[]� ^3�[]� �U��V��~ ��   W�}����   �$�؟�E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN�t��M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W��d  ���F    _^]� �� �.�<�O�^�m�|�����U��V��~ �  �E W�}�E����   �$�0����]������   �   ���]����A��   �   ���]����A��   �r���]������   �`�E������A��uN��������   �C�E��������u1������A{{�*�E���������E������A�����]����DzU����ءt��U�H0�F���   j j j j j j j RjP���E �U(��(R���\$�E�$W�c  ���F    _^]�$ �I *�?�T�f�x�������Ơ������������U���E �E�Uj���\$�E�\$�E�$PR�w���]�  ���U���E �E�Uj���\$�E�\$�E�$PR�G���]�  ���U���E �E�Uj���\$�E�\$�E�$PR����]�  ��̋�3�� <|�H�H�H�������������VW��3��<|9~u�t��H4�V�R�Ѓ��~�~_^����U��t��P4�E�I�RtPQ�҃�]� �U��U��t3�A�t��I0R���   P�ҋt��Q0�M���   QP�҃�]� �t��P0�E�I�R|PQ�҃�]� ������̡t��P4�A�JP�у������������̡t��P4�A�JP�у������������̡t��P4�A�JP�у������������̡t��P4�A�J|P�у������������̡t��P4�A���   P�у����������U��t��P4�E�I�RP�EP�EP�EPQ�҃�]� �����U��t��P4�E�I�RP�EP�EP�EPQ�҃�]� �����U��t��P4�E�I�R PQ�҃�]� �U��t��P4�E�I�R$PQ�҃�]� �U��t��P0�E�I���   P�EP�EP�EPQ�҃�]� ��U��t��P4�E�I���   PQ�҃�]� ��������������U��t��P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U��t��P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U��t��P4�E�I�R(PQ�҃�]� �U��t��P4�E�I�R,P�EP�EPQ�҃�]� ���������U��t��P4�E�I�R0P�EPQ�҃�]� ������������̡t��P4�A�J4P��Y��������������U����UV��EP�M�Q�NR�E�    �E�    �����t��H4�V�AR�Ћt��Q0�Rhj �M�Q�M�Q�M�Q�M�QP�F�HQ�҃� �} ^t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ��������������U��t��P4�E�I�R8PQ�҃�]� �U��t��P4�E�I�R<PQ�҃�]� �U��t��P4�E�I���   P�EPQ�҃�]� ����������U��t��E�P4�A��  ���$P�у�]� ��������̡t��P4�A�J@P�у������������̡t��P4�A��  P�у����������U��t��P4�E�I�RDP�EPQ�҃�]� �������������U��t��P4�E�I�RHP�EPQ�҃�]� �������������U��t��P4�E�I�RLP�EPQ�҃�]� �������������U��t��P4�E�I�RPP�EPQ�҃�]� �������������U��t�SV�uW�����   �QV�҃�����   �t����   �]�QS�҃�S��uA�t����   �Q@�ҋءt����   �Q@V�ҋt��Q4�JPSP�GP�у�_^[]� �t����   �H�у���uD�t����   �H8S�ыt��؋��   �H@V�ыt��J4�WSP�AHR�Ѓ�_^[]� hh|h�  ��   �t����   �BV�Ѓ�����   �t����   �]�BS�Ѓ�S��uC�t����   �B@�Ћt����   �؋B8V�Ћt��Q4�JLSP�GP�у�_^[]� �t����   �H�у���uD�t����   �H8S�ыt��؋��   �H8V�ыt��J4�WSP�ADR�Ѓ�_^[]� hh|h�  �
hh|h�  �t��Q��0  �Ѓ�_^[]� �U��t��P4�E�I��  P�EP�EP�EPQ�҃�]� ��U��t��P4�E,P�E(P�E$P�E �IP�E�RTP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U��t��P4�E�I�RXP�EP�EP�EPQ�҃�]� ����̡t��P4�A�J`P��Y�������������̡t��P4�A�JdP�у�������������U��t��P4�E�I��   P�EP�EP�EPQ�҃�]� ��U��t��P4�E�I�R\P�EP�EP�EP�EP�EPQ�҃�]� �������������U��t��P4�E�I�RhP�EPQ�҃�]� �������������U��t��P4�E�I��  P�EPQ�҃�]� ����������U��t��P4�E�I��  P�EPQ�҃�]� ����������U��t��P4�E�I�RpP�EPQ�҃�]� �������������U���,V��~ ��   �t��V�H4�AR�Ѓ} t �t��Q0�RlP�F�HQ�҃�^��]� ��hARDb�MԉE��E�    �\���P�M�Q�N�U�R�{����t����   ��U�R�Ѓ��M��m���^��]� ������U��t��P4�E�I�RlPQ�҃��   ]� ������������U��t��E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U��t��P4�E�I���   P�EP�EPQ�҃�]� �����̡t��P4�A���   P�у���������̸   ����������̸   �����������U��t�V��H4�V�A$h�  R�Ћt��Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U��t��P4�E�I�RxP�EP�EP�EPQ�҃�]� �����U��t��P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}�M���t�t��P���   j j���Љ�u��t�t��Q���   j j���Љ�t��Q4�E��H�RpVWQ�҃�_^[��]� �U��Q�t��P�B SVW�}���3���=INIb�/  �  =SACbvt+=$'  t
=MicM�  ��B$W����_�   ^��[��]� ��R3��E��E�EP�M�Q���҅�t�t��U�H4�E�R�VP�AR�Ѓ�_�   ^��[��]� =ARDb�  �t��Q���   j j���Ћt��Qj �؋��   j���Ћt��Qj �E����   j���Ћt��Qj �E���   j���ЋM���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>���I���P���!���P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� �t��Q���   j hIicM���ЋWP�B ����_^[��]� �������������U��t��P4�E�I�RTh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M��:����t��Q4�JlP�FP�у��M��\���^��]��������V����{�t��H0�Vh@o�҉F���F    ��|�F   ��^��������V��F��{��t�t��Q0P�B�Ѓ��F    ^������U��t��P�B VW�}�����=cksat`=ckhct�MQW��荽��_^]� �Nj j j j j j �F   �t��B0���   j j j Q�҃�(��t'_�F    �   ^]� �~ t��P����_^]� _3�^]� ���U��t��H���  ]��������������U��t��H0���   ]��������������U��t��H0�U�E��VWRP���   �U�R�Ћt��Q�u���BV�Ћt��Q�BVW�Ћt��Q�J�E�P�у�_��^��]������������U��t��H0���   ]��������������U��t��H0���   ]��������������U��t��H0���   ]��������������U��Ej0P�K  ��]��������������U��Ej0P�2�  ��P�iK  ��]�����U��E�M��j0PQ�U�R�7�  ��P�>K  �t��H�A�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P�c�  ��P��J  �t��Q�J�E�P�у���]��U��Ej$P��J  3Ƀ�������]����U��Ej$P�r�  ��P�J  3Ƀ�������]�����������U��E�M��Vj$PQ�U�R�f�  ��P�mJ  �t�3Ƀ��B�P����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P��  ��P�J  �t�3Ƀ��B�P����M�Q�҃���^��]����U��t��H�U�E���   RPj �у�]���������������U��t��H�U�ER�UP���   Rj �Ѓ�]�����������U��t��P4�E�I�R,P�EP�EPQ�҃�]� ���������U��t��P4�E�I�R0P�EPQ�҃�]� ������������̡t��P4�A�J4P��Y��������������U��U��V��EP�M�QR���4����t��H0�E�P� R�U�R�U�R�U�R�U�R�VP�AhR�Ѓ��} ^t(�} t(�E�M�;�~<�U��;�}3�E�M�;�~)�U���} u�E�M�;�~�U��;�}�   ��]� 3���]� �����������U��ESVW�؅�u�Y�t��P�}���   j hdiuM���Ћ���tK;3u	_^3�[]� �t��Q���   j hIicM����;�u�t��Q���   j h1icM���Шu��3_^�   []� �����U��t��P�BT��(V�uhfnic���Ѕ�t�t��Q�ȋ��   j
�Ѕ���   �t��Q�RPhfnic�E�P����P�M��ߴ���M�������u�E�P��������M������t��Q�B ���Ѓ��t�t��Q�B ���Ѕ�u�t��Q�B$hfnic���Ћt��E�Q�R8Pj
����^��]���������U��t��P0�E�IP�EP�EP�EPQ���   �у�]� ��U��t��P0�E�IV�p� ���   V�uj j j V�uVj Pj=Q�҃�(^]� ����U��t��P0�E�IV�p� ���   V�uV�uj j j�Vj Pj=Q�҃�(^]� ���̡t��I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V����{�t��H0�WVh@o�ҋ}�F�E�F    �F   ��|�F�t��Q���   ��j hmyal���ЉF��t��t�F    �t��Q���   j
hhfed���ЉF_��^]� �����������U��t��P�B VW�}�����=ytsdt�MQW�������_^]� �t��B0�N���   Q�ҋ�P������_�   ^]� ��3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ��������������������̸0}�����������U���E�Y(]� ���U���(V���P(�M�Q���ҋN��t&�t��R0j j j j j j P���   j jQ�Ѓ�(�t��Q�J�E�P�ыt��B�P�M�Q�ҋF����t �t��Q0�RHj �M�Qj jj?j P�҃��t��H�A�U�WR�Ћt��Q�J�E�P�ыF����u3��;�t��E�    �J0�U�Rj j j h  
 j�U�Rh�  jP���   �Ћ}���(�t��Q�J�E�P�у���_u3�^��]Ët��B�P�M�Q�ҋF����t �t��Q0�RHj �M�Qj j j8j P�҃��t��H�A�U�R�ЋF����t�t��Q0jP�BP�Ѓ��t��Q�J�E�P�у��M�詯��Ph   h  K j;�U�Rh	��h�  ���w����t��H�A�U�R�Ѓ��M��˯���F��t�t��Q0P�BX�Ѓ��F��t�t��Q0P�BX�Ѓ��F��t'�t��Q0j j j j j jj j jP���   �Ѓ�(j�v$�QA  ���   ^��]�����U���SV��W�~j���y�  ��V�^(3ۉ^4�^8�^<�t��H0�Ah�   R�Ћt��Q�J�E�P�ыt��B�PSj��M�h@}Q�҃�SS�E�P�M�Q���E��  �]��	����t��B�P�M�Q�҃�Sj����  _^[��]���̍A�������������U��VW��~4 tA�I �t��H��0  hh|hs  ��j
�oJ  �t��HP�V �AR�Ѓ���uQ9F4ut��QP�Bh�~0���Ѓ~4 t;�t��Q��0  hh|h�  �Ћt��QP�Bl�������m���_3�^]� �M�U�N8�V4�t��PP�Bl�~0���Ѓ~4 t%j
��I  �t��QP�F �JP�у���u�9F4uۋt��BP�PhS���ҋ^<�F<    �t��PP�Bl���Ћ�[_^]� ��U��t��P�B ��@VW�}�����=MicMtI=fnic��   j�M�������uP���=����M��%����t��Q�B4jj����_�   ^��]� �t��Q���   j hIicM����=�����   htats�M�蒬���t��Q�B0j j�M��ЍM�Q�U�R�E�P���E��  �E�    茳���t����   �
�E�P�у��M��}����F�F   ��t�t��J0�QP�҃��EPW���1���_^��]� ���������U��E��V��t3�^]� j�N�a�  j�
>  �F    �v����t�t��H0�QV�҃��   ^]� ��������������j����  j�=  ��3�����������U��E3�h�����h  ���P�Ej BR�Uj PR�����]� �U��Q�Q��u3���]� �E�H� V�5t�Q�M�Q�E�    �v0PR�V8�ҋ�����t@�E���t9�t��Q�M�RQP�ҋE�����t�t��QW��P�B��W�S  ��_��^��]� ������U��t���V��H�A�U�R�ЋU���M�QR���D�������u�t��H�A�U�R�Ѓ�3�^��]� �M�Q�M�����t��B�P�M�Q�҃���^��]� �������U��t���V��H�A�U�R�ЋU���M�QR��������M��t��P�R8�E�PQ�M�ҡt��H�A�U�R�Ѓ���^��]� �������������U���V��M��/����M�E�PQ��������t����B�U�@<�M�Q�MR�ЍM�������^��]� ����U��t��P�E���   Vj ��MP��h���h  �j j jj P�EP������^]� ��������������U��t�V�uW�����   �QV�҃�V��u,�t����   �Q@�ҋt��Q4�J P�GP�у�_^]� �t����   �H�у���u.�t����   �H8V�ыt��J4�WP�A$R�Ѓ�_^]� �t��Q��0  hh|h  �Ѓ�_^]� �����U���4�t��H�QSVW�}W�ҡt��P�u���   ��3�SS�Ή]�Ћt��QS�E����   j���Ћ�;��L  �d$ �} ~l�t��Q�J�E�P�ыt��B�Pj j��M�hD}Q�ҡt��P�B<�����Ћt��Q�RLj�j��M�QP���ҡt��H�A�U�R�Ѓ��t��Q0�E����   VP�M�Q�ҋ�t��H�A�U�R�Ћt��Q�J�E�PV�ыt��B�P�M�Q�ҡt��P�B<�����Ћt��Q�RLj�j��M�QP���ҡt��H�A�U�R�Ћt��Q�u���   �E��j ��
S���Ћt��Q���   �E�j �CP���ҋ����������_^[��]����������������U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj AQj R�UR������^]� ��������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR�ϯ��^]� ����������U��E�E43҃8��R�U<R�U(���\$�E,�$R�E �� �\$�E�\$�E�\$�@�E�$P�°��]�8 ��������������U��E�@3҃8��E��Rj ���T$�$htemf�E �� �\$�E�\$�E�\$�$P�g���]�  ���U��E�E 3҃8��R�� �\$�E�\$�E�\$�@�E�$P�
���]�  ������U��E�@3҃8��E��Rj ���T$�$htcpf�E �� ��v�����\$�E���\$�}�\$�$P�˯��]�  �������U��E3҃8��R�UR�UR�UR�UP�EPR����]� U��E3҃8V�u��V��RP�EP�����^]� ����������U��Q��u3�]� �E�E�H� V�5t��v0Q�M Q�M���\$���E�$QPR�V(�҃�$^]� ���U��t��P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U��t��P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U��t���P�E���   V���$��MP�ҋ���u�^�    ^]� ��u�^����D{�   ^]� ��^]� ������U���0��t��U�V�U���M�]��P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�Q�P�Q�P�@�Q�A����  ^��]� ��������U��� ��t��]�V���M�]��P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�@�Q�A����  ^��]� �����U���VW�}�M�;}us�t��P�u���   j htsem���Ѕ�uS�t��QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E��������t�E�M�P�w  _�   ^��]� _3�^��]� U���VW�}�M�;}us�t��P�u���   j htsem���Ѕ�uS�t��QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E�跲����t�E�M�P��  _�   ^��]� _3�^��]� U���SVW�}��;}uz�t��P�u���   j htsem���Ѕ�uZ�t��QP���   hrdem���Ѕ�u=��M�Q�]��M�U�R�}��E��e�����t�E������$�  _^�   [��]� _^3�[��]� ��������U���4�ESW�}�M�;�t;Et	;E��   �t��P�]���   j htsem���Ѕ���   �t��QP���   hrdem���Ѕ�uj�M��U�ỦE��UԉE��]܉E�M�E�P�M�Q�M�U�U�R�E�P�}��ѱ����t+�E̋M�������E��X�E��X��  �   _[��]� _3�[��]� ��������U���SVW�}��;}��   �t��P�u���   j htsem���Ѕ�uj�t��QP���   hrdem���Ѕ�uM��U�M��]���Q�M�]��E�R�E�P�}��H�����t%�E��������E��X�  �   _^[��]� _^3�[��]� ���̋A���X(Q�ȋB$��j j h���� 4  ���������������U��t���0VW���H�A�U�R�Ћt��Q�J�E�P�ыE���U�RP�M�Q�M�,B���t��J�U�RP�A�Ћt��Q�J�E�P�ыt��B�P�M�Q�ҡt��H�Q��V�ҡt��H�A�U�VR�Ѓ�����  �t��Q�J�E�P�у�_^��]� ������������U���SVW�}��;}��   �t��P�u���   j htsem���Ѕ�ue�t��QP���   hrdem���Ѕ�uH�t��Q�J�E�P�ыM���U�R�E�P�}��E�    �-�����u �t��Q�J�E�P�у�3�_^[��]� ���U��R�{@�����  �t��H�A�U�R�Ѓ�_^�   [��]� ��U��V�u���  ��^]� �����������U���L�t�SV��H�A�U�R�Ћt��Q�J3�Sj��E�hH}P���F(��v��S�U�SR�E��  �]��: P�E�P�T����P�M�Q�������P�U�R�������t��H�A�U�R�Ћt��Q�J�E�P�ыt��B�P�M�Q�҃�htats�M��=����t��P�B0jj�M����F(�t��Q�B,���$j�M��ЍM�Q�U�R�E�P���E��  �]�� ����t����   �
�E�P�у�9^4t^�t��BP�PhW�~0���ҋF4;�t�N8Q�Ѓ��F<�^8�^4��t��B��0  hh|h�  �у��t��BP�Pl����_�M�讛��^[��]� ������U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�E�Y����D{�   ]� �����������U�����u�E�    �Y�E�Y�E�Y]� ��u-�E�Y����Dz�E�Y����Dz�E�Y����D{�   ]� �����U��V�����u#�E�M�U�F�E�N�V�    �F^]� ��u�MQ�VR�O�������t�   ^]� �������������U��V��~ �<|u�t��H4�V�R�Ѓ��E�F    �F    t	V�q  ����^]� �������U��V��F��{��t�t��Q0P�B�Ѓ��E�F    t	V�(  ����^]� ��������������U���V��3ɍF��H������t��M��M����   �RQ�M�QP�ҡt����   ��U�R�Ѓ���^��]��������������U��V�����u �    �t��H�A���UVR�Ѓ��#��u�t��Q�Rx�EP�N�҅�t�   �t��H�A�UR�Ѓ�^]� �������U��V�u���t�t��QP��Ѓ��    ^]���������̡t��H��@  hﾭ���Y����������U��E��t�t��QP��@  �Ѓ�]����������������U��t��H���  ]��������������U��t��H��  ]�������������̡t��H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�6 ������u_^]Ã} tWj V� ��_������F�x�   ^]���U��t��E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�5 ������u_^]�Wj V� ��_������F�x�   ^]�������������U��t��E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�5 ������u_^]�Wj V�& ��_������F�x�   ^]�������������U��t��E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�4 ������u_^]�Wj V� ��_������F�x�   ^]�������������U��t��E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�4 ������u_^]�Wj V�& ��_������F�x�   ^]�������������U��M��t-�=x� t�y���A�uP�A ��]át��P�Q�Ѓ�]��������U��M��t-�=x� t�y���A�uP� ��]át��P�Q�Ѓ�]��������U��t��H�U�R�Ѓ�]���������U��t��H�U�R�Ѓ�]���������U��t��E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��2 ������u_^]�Wj V�� ��_������F�x�   ^]���������U��t��E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   �t���t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��1 ������u_^]�Wj V�� ��_������F�x�   ^]����������U��E��w�   �t���t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�P1 ������u_^]�Wj V�` ��_������F�x�   ^]�������U��t��H�U�R�Ѓ�]���������U��t��H�U�R�Ѓ�]���������U��t��H�U�R�Ѓ�]���������U��t��H�U�R�Ѓ�]��������̡t��HL���   ��U��t��H@�AV�u�R�Ѓ��    ^]�������������̡t��HL�������U��t��H@�AV�u�R�Ѓ��    ^]�������������̡t��PL���   Q�Ѓ�������������U��t��PL�EP�EPQ���   �у�]� �������������U��t�V��HL���   V�҃���u�t��U�HL���   j RV�Ѓ�^]� �t����   �ȋBP�Ћt����   �MP�BH��^]� �����̡t��PL��(  Q�Ѓ�������������U��t��PL�EP�EPQ��,  �у�]� ������������̡t��HL�Q�����U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��PL�E�R��VPQ�M�Q�ҋu��P���e����M��}�����^��]� ����U��t��PL�EPQ���   �у�]� �U��t��PL�EP�EPQ�J�у�]� �t��PL�BQ�Ѓ���������������̡t��PL�BQ�Ѓ���������������̡t��PL�BQ�Ѓ����������������U��t��PL�EP�EP�EPQ�J �у�]� ������������U��t��PL�EPQ��4  �у�]� �U��t��PL�EP�EP�EPQ�J$�у�]� ������������U��t��PL�EP�EP�EP�EPQ�J(�у�]� �������̡t��PL�B,Q�Ѓ���������������̡t��PL�B0Q�Ѓ����������������U��t��PL�EP�EPQ��  �у�]� ������������̡t��PL���   Q�Ѓ�������������U��t��PL�E��  ��VPQ�M�Q�ҋu��P���B����M��Z�����^��]� ̡t��PL�B4Q�Ѓ���������������̡t��PL�B8j Q�Ѓ��������������U��t��PL���   ]��������������U��t��PL���   ]��������������U��t��PL���   ]��������������U��t��PL���   ]��������������U��t��PL���   ]��������������U��t��PL���   ]��������������U��t��PL��l  ]��������������U��t��PL���   ]��������������U��t��PL���   ]��������������U��t��PL���   ]��������������U��t��PL�EPQ�J<�у�]� ���̡t��PL�BQ��Y�U��t��PL�EP�EPQ�J@�у�]� U��t��PL�Ej PQ�JD�у�]� ��U��t��PL�Ej PQ�JH�у�]� ��U��t��PL�EjPQ�JD�у�]� ��U��t��PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��E  W�M�Q�U�R���tM  ���M����7  ��t�t����   ��U�R�Ѓ�_^3�[��]Ët����   �J8�E�P�ыt������   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  ��D  j�M�Q�U�R����L  �M���6  �t����   ��U�R�Ѓ�^��]�����������U���$�t��UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��zD  j�E�P�M�Q���YL  �M��q6  �t����   ��M�Q�҃�_^��]� ��U���$�t��UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}���C  j�E�P�M�Q����K  �M���5  �t����   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��C  W�M�Q�U�R���TK  ���M����5  ��t+�u���f���t����   ��U�R�Ѓ�_��^[��]� �t����   �JL�E�P�ыu��P���%g���t����   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}���B  W�M�Q�U�R���J  ���M�����4  ��t+�u����e���t����   ��U�R�Ѓ�_��^[��]� �t����   �JL�E�P�ыu��P���ef���t����   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��B  W�M�Q�U�R����I  ���M����4  _^��[t�t����   ��U�R�������]Ët����   �J<�E�P���]��t����   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��dA  W�M�Q�U�R���$I  ���M����W3  ��t�t����   ��U�R�Ѓ�_^3�[��]Ët����   �J8�E�P�ыt������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��@  W�M�Q�U�R���tH  ���M����2  ��t-��u�t�����   ���^�U�R�Ѓ�_��^[��]� �t����   �JP�E�P�ы�u�H��P�@�N�t��V���   �
�F�E�P�у�_��^[��]� �����̡t��PL���   Q��Y��������������U��t��PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U��t��PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��$?  W�M�Q�U�R����F  ���M����1  ��t-��u�t�����   ���^�U�R�Ѓ�_��^[��]� �t����   �JP�E�P�ы�u�H��P�@�N�t��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��T>  W�M�Q�U�R���F  ���M����G0  ��t-��u�t�����   ���^�U�R�Ѓ�_��^[��]� �t����   �JP�E�P�ы�u�H��P�@�N�t��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��=  W�M�Q�U�R���DE  ���M����w/  ��t-��u�t�����   ���^�U�R�Ѓ�_��^[��]� �t����   �JP�E�P�ы�u�H��P�@�N�t��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��<  W�M�Q�U�R���tD  ���M����.  ��t�t����   ��U�R�Ѓ�_^3�[��]Ët����   �J8�E�P�ыt������   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  ��;  j�M�Q�UR����C  �M��-  �t����   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��;  j�U�R�E�P���nC  �M��-  �t����   �
�E�P�у�^��]� ��������U���$�t��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
;  j�E�P�M�Q����B  �M��-  �t����   ��M�Q�҃�_^��]� ��U���$�t��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��:  j�E�P�M�Q���iB  �M��,  �t����   ��M�Q�҃�_^��]� ��U���$�t��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
:  j�E�P�M�Q����A  �M��,  �t����   ��M�Q�҃�_^��]� ��U���$�t��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��9  j�E�P�M�Q���iA  �M��+  �t����   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��9  j�U�R�E�P����@  �M��+  �t����   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}��8  W�M�Q�U�R���t@  ���M����*  ��t-��u�t�����   ���^�U�R�Ѓ�_��^[��]� �t����   �JP�E�P�ы�u�H��P�@�N�t��V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���7  W�M�Q�U�R���?  ���M�����)  ��t�t����   ��U�R�Ѓ�_^3�[��]Ët����   �J8�E�P�ыt������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��47  W�M�Q�U�R����>  ���M����')  ��t�t����   ��U�R�Ѓ�_^3�[��]Ët����   �J8�E�P�ыt������   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ���̡t��PL���  ��U���$�t��UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��:6  j�E�P�M�Q���>  �M��1(  �t����   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���5  j�U�R�E�P���=  �M���'  �t����   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��_5  j�U�R�E�P���>=  �M��V'  �t����   �
�E�P�у�^��]� ��������U��t��H���   ]��������������U��t��H���   ]�������������̡t��H���   ��t��H���   ��U��t��H���   V�u�R�Ѓ��    ^]�����������U��t��H���   ]��������������U��t��HL�QV�ҋ���u^]át��H�U�Ej R�UP��h  RV�Ѓ���u�t��Q@�BV�Ѓ�3���^]��������U��t��H�U�E��h  j R�U�� P�ERP�у�]����U��t��H���   ]��������������U��t��H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡t��PL�BLQ�Ѓ���������������̡t��PL�BPQ�Ѓ����������������U��t��PL�EP�EPQ�JT�у�]� U��t��PL�EPQ��  �у�]� �U��t��PL�EPQ���   �у�]� ̡t��PL�BXQ�Ѓ����������������U��t��PL�EP�EP�EPQ�J\�у�]� ������������U���4�t�SV��HL�QW�ҋ�3ۉ}�;��x  �M��!x���t��E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡt����   �BSSW���Ѕ���   �t��QL�BW�Ћ���;���   ��    �t����   �B(���ЍM�Qh�   ���u��j  ������   �M�;���   �t����   ���   S��;�tm�t����   �ȋB<V�Ћt����   ���   �E�P�у�;�t�t��B@�HV�у���;��\����}��M��!  �M��Yw����_^[��]� �}��t��B@�HW�ыt����   ���   �M�Q�҃��M��9!  �M��w��_^3�[��]� �����̡t��PL�B`Q�Ѓ���������������̡t��PL�BdQ�Ѓ����������������U��t��PL�EPQ�Jh�у�]� ���̡t��PL��D  Q�Ѓ������������̡t��PL�BlQ�Ѓ����������������U��t��PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh �h �h��h��R�Q�U R�UR�UR�U���A�$�5t��vLRP���   Q�Ѓ�4^]�  ������̡t��PL���   Q�Ѓ�������������U��t��PL�EP�EP�EPQ��   �у�]� ���������U��t��PL��H  ]�������������̡t��PL��L  ��U��t��PL��P  ]��������������U��t��PL��T  ]��������������U��t��PL��p  ]��������������U��t��PL��t  ]��������������U��t��PL�EP�EP�EP�EP�EPQ���   �у�]� �U��t��PL�EP�EP�EPQ���   �у�]� ���������U��t��PL�EP�EP�EP�EPQ��   �у�]� �����U��t��HL���   ]��������������U��t��HL���   ]��������������U��t��HL���   ]�������������̡t��HL��  ��t��HL��@  ��U��t��PL���  ]��������������U��t��PL���  ]��������������U��t��PL���  ]��������������U��� �t�V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\�t��QLjP���   ���ЋM��U�Rh=���M�}��  ���t����   ���   �U�R�Ѓ��M��u��  ��_^��]Ët����   ���   �E�P�у��M��u��^  _�   ^��]����U��� �t�V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\�t��QLjP���   ���ЋM��U�Rh<���M�}��C  ���t����   ���   �U�R�Ѓ��M��u��  ��_^��]Ët����   ���   �E�P�у��M��u��  _�   ^��]����U��t��P8�EPQ�JD�у�]� ���̡t��H8�Q<�����U��t��H8�A@V�u�R�Ѓ��    ^]�������������̡t��H8�������U��t��H8�AV�u�R�Ѓ��    ^]��������������U��t��P8�EP�EP�EPQ�J�у�]� ������������U��t��P8�EP�EPQ�J�у�]� �t��P8�BQ�Ѓ����������������U��t��P8�EPQ�J �у�]� ����U��t��P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U��t��P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U��t��P8�EP�EPQ�J(�у�]� U��t��P8�EP�EP�EPQ�J,�у�]� ������������U��t��P8�EP�EP�EPQ�J�у�]� ������������U��t��P8�EP�EP�EP�EP�EPQ�J�у�]� ����U��t��P8�EP�EPQ�J0�у�]� U��t��P8�EP�EP�EPQ�J4�у�]� ������������U��t��P8�EPQ�J8�у�]� ����U��t��H��x  ]��������������U��t��H��|  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H�A,]�����������������U��t��H���  ]��������������U��t��H�QV�uV�ҡt��H�Q8V�҃���^]�����̡t��H�Q<�����U��t��H�I@]����������������̡t��H�QD����̡t��H�QH�����U��t��H�AL]�����������������U��t��H�IP]�����������������U��t��H��<  ]��������������U��t��H��,  ]��������������U��t��H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡t��H���   ��t��H���  ��U��t��H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U��t��H�A]�����������������U��t��H��\  ]��������������U��t��H�AT]�����������������U��t��H�AX]�����������������U��t��H�A\]����������������̡t��H�Q`�����U��t��H���  ]�������������̡t��H�Qd����̡t��H�Qh�����U��t��H�Al]�����������������U��t��H�Ap]�����������������U��t��H�At]�����������������U��t��H��D  ]��������������U��t��H��  ]��������������U��t��H�Ix]�����������������U��t��H��@  ]��������������U��V�u���G���t��H�U�A|VR�Ѓ���^]���������U��t��H���   ]��������������U��t��H��h  ]��������������U��t��H��d  ]��������������U��t��H���  ]�������������̡t��H���   ��U��t��H��l  ]��������������U��t��H��   ]��������������U��t��H��  ]��������������U��V�u����h���t��H���   V�҃���^]���������̡t��H��`  ��U��t��H��  ]��������������U��t��H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U��t��H���  ]��������������U��U�E�t��H�E���   R���\$�E�$P�у�]�U��t��H���   ]��������������U��t��H���   ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���   ]��������������U��t��H���   ]��������������U��t��H���   ]��������������U��t��H���   ]��������������U��t��H���   ]��������������U��t��H���   ]��������������U��t��P���E�P�E�P�E�PQ���   �у����#E���]����������������U��t��P���E�P�E�P�E�PQ���   �у����#E���]����������������U��t��P���E�P�E�P�E�PQ���   �у����#E���]����������������U��t��H��8  ]��������������U��V�u(V�u$�E�@�t��R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@�t��R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��t��P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U��t��P0�EP�EP�EP�EPQ���   �у�]� ����̡t��P0���   Q�Ѓ�������������U��t��P0�EP�EPQ���   �у�]� �������������U��t��P0�EP�EP�EP�EPQ���   �у�]� ����̡t��P0���   Q�Ѓ������������̡t��H0���   ��U��t��H0���   V�u�R�Ѓ��    ^]�����������U��t��H��H  ]��������������U��t��H��T  ]�������������̡t��H��p  ��t��H���  ��U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H�U�E��X  ��VR�UPR�E�P�ыu�    �F    �t����   �Qj PV�ҡt����   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M��Jb��P�E�hicMCP�k������M��pb���t����   �JT�E�P�у���u(�u����a���t����   ��M�Q�҃���^��]át����   �AT�U�R�Ћu��P����a���t����   �
�E�P�у���^��]�������������U��t��H��  ]��������������U��t��H��\  ]��������������U��t��H�U��t  ��V�uVR�E�P�у����S@���M��?����^��]�����U��t��H�U���  ��VWR�E�P�ыt��u���B�HV�ыt��B�HVW�ыt��B�P�M�Q�҃�_��^��]����������������U��t��H�U���  ��VWR�E�P�ыt��u���B�HV�ыt��B�HVW�ыt��B�P�M�Q�҃�_��^��]����������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H�U�E��VWj R�UP�ERP��t  �U�R�Ћt��Q�u���BV�Ћt��Q�BVW�Ћt��Q�J�E�P�у�(_��^��]��U��t��H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    �t����   j P�BV�Ћt����   �
�E�P�у�$��^��]���U��t��H��8  ]��������������U���  ��3ŉE��M�EPQ������h   R�� ����|	=�  |#��t��H��0  hP}hH  �҃��E� �t��H��4  ������Rh�}�ЋM�3̓���  ��]�������U��t��H��  ��V�U�WR�Ћt��Q�u���BV�Ћt��Q�BVW�Ћt��Q�J�E�P�у�_��^��]����U��t��H��  ��V�U�WR�Ћt��Q�u���BV�Ћt��Q�BVW�Ћt��Q�J�E�P�у�_��^��]����U��t��H��p  ��$�҅�trh���M��)]���t��P�E�R4Ph���M��ҡt��P�E�R4Ph���M���j �E�P�M�hicMCQ�����t����   ��M�Q�҃��M��]����]�U��t��H��p  ��$V�҅�u�t��H�u�QV�҃���^��]�Wh!���M��|\���t��P�E�R4Ph!���M���j �E�P�M�hicMCQ�����t����   �QHP�ҋu���t��H�QV�ҡt��H�QVW�ҡt����   ��U�R�Ѓ�$�M��=\��_��^��]������U��t��H��p  ��$V�҅�u�t��H�u�QV�҃���^��]�Wh����M��[���t��P�E�R4Ph����M���j �E�P�M�hicMCQ�����t����   �QHP�ҋu���t��H�QV�ҡt��H�QVW�ҡt����   ��U�R�Ѓ�$�M��m[��_��^��]������U��t��H��p  ��$�҅�u��]�Vh#���M���Z���t��P�E�R4Ph#���M���j �E�P�M�hicMCQ������t����   �Q8P�ҋ�t����   ��U�R�Ѓ��M���Z����^��]���������������U��t��H��p  ��$�҅�u��]�Vhs���M��TZ���t��P�E�R4Phs���M���j �E�P�M�hicMCQ�W����t����   �Q8P�ҋ�t����   ��U�R�Ѓ��M��5Z����^��]���������������U��t��H���  ]��������������U��t��H��@  ]��������������U��t��H���  ]��������������U��V�u���t�t��QP��D  �Ѓ��    ^]������U��t��H��H  ]��������������U��t��H��L  ]��������������U��t��H��P  ]��������������U��t��H��T  ]��������������U��t��H��X  ]��������������U��t��H��\  ]�������������̡t��H��d  ��U��t��H��h  ]��������������U��t��H��l  ]�������������̡t��H���  ��U��t��H�U���  ��VR�E�P�ыu��P���#X���M��;X����^��]�����U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H��l  ]��������������U��t��H���  ]��������������U��t��H���  ]��������������U��t��H��$  ]��������������U��t��H��(  ]��������������U��t��H��,  ]�������������̡t��H��0  ��t��H��<  ��U��t��H���  ]�������������̡t��H���  ��U��t��H���  ]������������������������������U��t��H��  ]�������������̡t��H��P  ��U��t��H��`  ]�������������̡t����   ���   ��Q��Y��������U��t��H�A�U��� R�Ћt��Q�Jj j��E�h�}P�ыUR�E�P�M�Q�m���t��B�P�M�Q�ҡt��H�A�U�R�Ћt��Q�J�E�P�у�,��]��h|�PhD ���  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h|�jhD ��  ����t
�@��t]��3�]��������Vh|�j\hD ���  ����t�@\��tV�Ѓ���^�����Vh|�j`hD ���  ����t�@`��tV�Ѓ�^�������U��Vh|�jdhD ���Y  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh|�jhhD ���  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh|�jlhD ����~  ����t�@l��tV�Ѓ�^�������U��Vh|�h�   hD ���~  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh|�h�   hD ���V~  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh|�jphD ���	~  ����t�@p��t�MQV�Ѓ�^]� ���^]� ��U��Vh|�jxhD ����}  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh|�j|hD ���}  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh|�j|hD ���I}  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� �������������U���Vh|�h�   hD ����|  ����t=���   ��t3�MQ�U�VR��h|�j`hD ��|  ����t�@`��t	�M�Q�Ѓ���^��]� �����̋���������������h|�jhD �|  ����t	�@��t��3��������������U��V�u�> t+h|�jhD �C|  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h|�jhD �|  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh|�jhD ���{  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh|�jhD ���y{  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh|�j hD ���<{  ����t�@ ��tV�Ѓ�^�3�^���Vh|�j$hD ���{  ����t�@$��tV�Ѓ�^�3�^���U��Vh|�j(hD ����z  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh|�j,hD ���z  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh|�j(hD ���Iz  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh|�j4hD ����y  ����t�@4��tV�Ѓ�^�3�^���U��Vh|�j8hD ����y  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh|�j<hD ���yy  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh|�jDhD ���<y  ����t�@D��tV�Ѓ�^�3�^���U��Vh|�jHhD ���	y  ����t�M�PHQV�҃�^]� U��Vh|�jLhD ����x  ����u^]� �M�PLQV�҃�^]� �����������U��Vh|�jPhD ���x  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh|�jThD ���\x  ����u^Ë@TV�Ѓ�^���������U��Vh|�jXhD ���)x  ����t�M�PXQV�҃�^]� U��Vh|�h�   hD ����w  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh|�h�   hD ���w  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh|�h�   hD ���Vw  ����u^]� �M���   QV�҃�^]� �����U��Vh|�h�   hD ���w  ����u^]� �M���   QV�҃�^]� �����U��Vh|�h�   hD ����v  ����u^]� �M���   QV�҃�^]� �����U��Vh|�h�   hD ���v  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh|�h�   hD �Uv  ����u�t��H�u�QV�҃���^��]ËM���   WQ�U�R�Ћt��Q�u���BV�Ћt��Q�BVW�Ћt��Q�J�E�P�у�_��^��]��U��Vh|�h�   hD ����u  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh|�h�   hD ���vu  ����t���   ��t�MQ����^]� 3�^]� �U��Vh|�h�   hD ���6u  ����t���   ��t�MQ����^]� 3�^]� �U��Vh|�h�   hD ����t  ����t���   ��t�MQ����^]� 3�^]� �Vh|�h�   hD ���t  ����t���   ��t��^��3�^����������������U��Vh|�h�   hD ���vt  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh|�h�   hD ���&t  ����t���   ��t�MQ����^]� ��������U��Vh|�h�   hD ����s  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh|�h�   hD ���s  ����t���   ��t��^��3�^����������������VW��3����$    �h|�jphD �Os  ����t�@p��t	VW�Ѓ������8 tF��_��^�������U��SW��3�V��    h|�jphD ��r  ����t�@p��t	WS�Ѓ������8 tqh|�jphD ��r  ����t�@p��t�MWQ�Ѓ�������h|�jphD �r  ����t�@p��t	WS�Ѓ�����V���������tG�]����E^��t�8��~=h|�jphD �Nr  ����t�@p��t	WS�Ѓ������8 u_�   []� _3�[]� ����������U��Vh|�j\hD ����q  ����t3�@\��t,V��h|�jxhD ��q  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh|�j\hD ���q  ����t3�@\��t,V��h|�jdhD �wq  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh|�j\hD ���6q  ����tG�@\��t@V�ЋEh|�jdhD �E��E�    �E�    � q  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh|�j\hD ���p  ����t\�@\��tUV��h|�jdhD �p  ����t�@d��t
�MQV�Ѓ�h|�jhhD �np  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh|�j\hD ���)p  ������   �@\��t~V��h|�jdhD �p  ����t�@d��t
�MQV�Ѓ�h|�jhhD ��o  ����t�@h��t
�URV�Ѓ�h|�jhhD �o  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh|�jthD ���vo  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h|�j`hD �>o  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh�����_�����^��]� ������U���Vh|�h�   hD ��n  ����tU���   ��tK�M�UQR�M�Q�Ћu��P������h|�j`hD �n  ����t%�@`��t�U�R�Ѓ���^��]ËE�uP���k�����^��]�����U���Vh|�h�   hD ���Sn  ����tR���   ��tH�MQ�U�R���ЋuP������h|�j`hD �n  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    �'�����^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t�t����   P�B@��]� �E��t�t����   P�BD��]� �t����   R�PD��]� �����U��t��P@�Rd]�����������������U��t��P@�Rh]�����������������U��t��P@�Rl]�����������������U��t��P@�Rp]�����������������U��t����   ���   ]�����������U��t����   ���   ]����������̡t��P@�Bt����̡t��P@�Bx�����U��t��P@�R|]����������������̡t��P@���   ��t����   �Bt��U��t��P@���   ]�������������̡t��P@���   ��U��t��P@���   ]��������������U��t��P@���   ]��������������U��t��P@���   ]��������������U��t��P@���   ]��������������U��t��P@���   ]��������������U��t��P@���   ]��������������U��t�V��H@�QV�ҋM����t��#����t��Q@P�BV�Ѓ�^]� �̡t��PH���   Q�Ѓ�������������U��t��P@�EPQ�JL�у�]� ���̡t��P@�BHQ�Ѓ����������������U��t��P@�EP�EP�EPQ�J�у�]� ������������U��t��P@�EPQ�J�у�]� ����U��t��P@�EP�EPQ�J�у�]� U��t��P@�EPQ�J �у�]� ����U��t����   �R]��������������U��t����   �R]��������������U��t����   �R ]��������������U��t����   ���   ]�����������U��t����   ��D  ]�����������U��t��E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U��t����   ���   ]����������̡t����   �B$��t��H@�Q0�����U��t��H@�A4j�URj �Ѓ�]����U��t��H@�A4j�URh   @�Ѓ�]�U��t��H@�U�E�I4RPj �у�]�̡t��H|�������U��V�u���t�t��Q|P�B�Ѓ��    ^]��������̡t��H|�Q �����U��V�u���t�t��Q|P�B(�Ѓ��    ^]��������̡t��H@�Q0�����U��V�u���t�t��Q@P�B�Ѓ��    ^]���������U��t��H@���   ]��������������U��V�u���t�t��Q@P�B�Ѓ��    ^]��������̡t��PH���   Q�Ѓ�������������U��t��PH�EPQ��d  �у�]� �U��t��H �IH]�����������������U��}qF uHV�u��t?�t����   �BDW�}W���Ћt��Q@�B,W�Ћt��Q�M�Rp��VQ����_^]����������̡t��P@�BT�����U��t��P@�RX]�����������������U��t��P@�R\]����������������̡t��P@�B`�����U��t��H��T  ]��������������U��t��H@�U�A,SVWR�Ћt��Q@�J,���EP�ыt��Z��h��hE  �΋��v;��Ph��hE  ���d;��P��T  �Ѓ�_^[]����U��t��PT�EP�EPQ�J�у�]� U��t��PT�EPQ�J�у�]� ����U��t��PT�EPQ�J�у�]� ����U��t��PT�E�R<��PQ�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��t��HT�]��U��t��H@�AV�u�R�Ѓ��    ^]�������������̡t��HT�hG  �҃�������������U��t��H@�AV�u�R�Ѓ��    ^]�������������̡t��PD�BQ�Ѓ���������������̡t��PD�BQ�Ѓ���������������̡t��PD�BQ�Ѓ����������������U��t��PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U��t��PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��t��PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��t��PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U��t��PX�EPQ�J�у�]� ����U��t��PX�EPQ�J�у�]� ����U��t��PX�EPQ�J�у�]� ����U��t��PX�EPQ�J�у�]� ����U��t��PX�EPQ�J$�у�]� ����U��t��PX�EPQ�J �у�]� ����U��t��PD�EP�EPQ�J�у�]� U��t��HD�U�j R�Ѓ�]�������U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��HD�	]��U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��HD�U�j R�Ѓ�]�������U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��U�HD�Rh2  �Ѓ�]����U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��U�HD�RhO  �Ѓ�]����U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��U�HD�Rh'  �Ѓ�]����U��t��H@�AV�u�R�Ѓ��    ^]�������������̡t��HD�j h�  �҃�����������U��t��H@�AV�u�R�Ѓ��    ^]�������������̡t��HD�j h:  �҃�����������U��t��H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E��t����   �R�E�Pj�����#E���]�̡t��HD�j h�F �҃�����������U��t��H@�AV�u�R�Ѓ��    ^]�������������̡t��HD�j h�_ �҃�����������U��t��H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E��t��E�    ���   �R�E�Pj������؋�]� ̡t��PD�B$Q�Ѓ���������������̡t��PD�B(Q�Ѓ���������������̡t��PD�BQ�Ѓ���������������̡t��PD�B(Q�Ѓ���������������̡t��PD�BQ�Ѓ���������������̡t��PD�B(Q�Ѓ���������������̡t��PD�BQ�Ѓ���������������̡t��PD�B(Q�Ѓ���������������̡t��PD�BQ�Ѓ���������������̡t��PD�B(Q�Ѓ���������������̡t��PD�BQ�Ѓ���������������̡t��PD�B(Q�Ѓ���������������̡t��PD�BQ�Ѓ���������������̡t��PD�B(Q�Ѓ���������������̡t��PD�BQ�Ѓ���������������̡t��PD�B(Q�Ѓ���������������̡t��PD�BQ�Ѓ���������������̡t��PD�B(Q�Ѓ���������������̡t��PD�BQ�Ѓ����������������U��t��H �Ah]�����������������U��t��H@�AV�u�R�Ѓ��    ^]�������������̡t��H �������U��V�u���t�t��Q P�B�Ѓ��    ^]���������U��t��P �EPQ�J4�у�]� ����U��t��P �EPQ�J�у�]� ����U��t��P �EPQ�J�у�]� ���̡t��P �BQ��Y�U��V�uW�����//���t��H �QVW�҃�_��^]� �����U��t��P �EPQ�J �у�]� ���̡t��P �B,Q�Ѓ���������������̡t��P �B0Q�Ѓ���������������̡t��H\�������U��t��H\�AV�u�R�Ѓ��    ^]�������������̡t��P\�BQ�Ѓ���������������̡t��P\�BQ�Ѓ����������������U��t��P\�EPQ�J�у�]� ����U��t��P\�EP�EPQ�J�у�]� U��t��P\�EPQ�J�у�]� ���̡t��P\�BQ�Ѓ����������������U��t��P\�EPQ�J �у�]� ����U��t��P\�EP�EPQ�J$�у�]� U��t��P\�EP�EP�EPQ�J(�у�]� ������������U��t��P\�EPQ�J0�у�]� ����U��t��P\�EPQ�J@�у�]� ����U��t��P\�EPQ�JD�у�]� ����U��t��P\�EPQ�JH�у�]� ���̡t��P\�B4Q�Ѓ����������������U��t��P\�EP�EPQ�J8�у�]� U��t��P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu���$���t��H\�QV�҃���S���$��3���~=��I �t��H\�U�R�U��EP�A(VR�ЋM��Q���$���U�R���}$��F;�|�_^[��]� ���������������U���VW�}�E��P��� ���}� ��   �t��Q\�BV�Ѓ��M�Q��� ���E���t]S3ۅ�~H�I �UR���e ���E�P���Z ���E;E�!���t��Q\P�BV�ЋE@��;E��E~�C;]�|�[_�   ^��]� _�   ^��]� U��t��E�PH�B���$Q�Ѓ�]� ���������������U��t��PH�EPQ���   �у�]� �U��t��PH�EPQ���  �у�]� �U��t��PH�EPQ���  �у�]� �U��t��PH�EP�EPQ��  �у�]� �������������U��t��PH�EP�EPQ��  �у�]� ������������̡t��PH���  Q�Ѓ�������������U��t��PH�EPQ���  �у�]� ̡t��PH���   j Q�Ѓ�����������U��t��PH�EPj Q���   �у�]� ��������������̡t��PH���   jQ�Ѓ�����������U��t��PH�EPjQ���   �у�]� ��������������̡t��PH���   jQ�Ѓ����������U��t��PH�EPjQ���   �у�]� ���������������U��t��PH�EP�EPQ���   �у�]� �������������U��t��PH�EP�EPQ���   �у�]� ������������̡t��PH���   Q�Ѓ�������������U��t��PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP��� ���������t�E�t��QH���   PVW�у���_^]� �����U��EVW���MPQ�,���������t�M�t��BH���   QVW�҃���_^]� ̡t��PH���   Q�Ѓ������������̡t��PH���   Q�Ѓ�������������U��t��PH�EPQ���   �у�]� �U��t��PH�EPQ���   �у�]� �U��t��PH�EP�EPQ��8  �у�]� �������������U��t��PH�EP�EPQ��   �у�]� ������������̡t��PH���  Q�Ѓ������������̡t��PH���  Q�Ѓ������������̡t��PH���  Q�Ѓ������������̡t��PH��  Q�Ѓ������������̡t��PH��  Q�Ѓ�������������U��t��PH�EP�EPQ��  �у�]� �������������U��t��PH�EP�EP�EPQ��   �у�]� ���������U��t��PH�EP�EP�EP�EPQ��|  �у�]� �����U��t��PH�EPQ��  �у�]� ̡t��PH��T  Q�Ѓ�������������U��t��PH�EP�EPQ��  �у�]� �������������U��t��PH�EPQ��8  �у�]� �U��t��PH�EPQ��<  �у�]� �U��t��PH�EP�EP�EPQ��@  �у�]� ���������U��t��PH�EPQ���  �у�]� ̡t��PH��L  Q��Y��������������U��t��PH�EPQ��H  �у�]� ̡t�V��H@�Q,WV�ҋt��Q��j �ȋ��   h�  �Ћt��QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡t��P@�B,Q�Ћt��Q��j �ȋ��   h�  �������U��t��E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��t��E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��t��PH�EP�EP�EPQ��   �у�]� ��������̡t��HH��  ��U��t��HH��  ]��������������U��t��E�PH��$  ���$Q�Ѓ�]� �����������̡t��PH��(  Q�Ѓ�������������U��t��PH�EP�EPQ��,  �у�]� �������������U��t��E�PH�EP�E���$PQ��0  �у�]� ���̡t��PH���  Q�Ѓ������������̡t��PH��4  Q�Ѓ������������̋��     �������̡t��PH���|  jP�у���������U��t��UV��HH��x  R��3Ƀ������^��]� ��̡t��PH���|  j P�у��������̡t��PH��P  Q�Ѓ������������̡t��PH��T  Q�Ѓ������������̡t��PH��X  Q�Ѓ�������������U��t��PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡t��PH��`  Q�Ѓ�������������U��t��PH�EPQ��d  �у�]� �U��t��E�PH��h  ���$Q�Ѓ�]� ������������U��t��E�PH��t  ���$Q�Ѓ�]� ������������U��t��E�PH��l  ���$Q�Ѓ�]� ������������U��t��PH�EPQ��p  �у�]� �U��t��PH�EP�EP�EP�EPQ���  �у�]� �����U��t��PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U��t��E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E�t��HH�E���   R�U���$P�ERP�у�]����������������U���E�M��}�<�  �M;�|�M;�~��]�����������U��t��PH�E���   Q�MPQ�҃�]� ������������̡t��PH���   Q��Y�������������̡t��PH���   Q�Ѓ������������̡t��PH���   Q��Y��������������U��t��PH�EP�EPQ���   �у�]� �������������U��t��PH�EP�EP�EP�EP�EPQ���  �у�]� ̡t��PH��t  Q��Y�������������̋�� �}�@    ���}�t��Pl�A�JP��Y��������U��t�V��Hl�V�AR�ЋE����u
�   ^]� �t��Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uËt��QlP�B�Ѓ�������U��t��Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E�t��HH�ER�U���$P���  R�Ѓ�]����U��t��HH���  ]��������������U��t��HH���  ]��������������U��U0�E(�t��HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U��t��HH���  ]��������������U��t��E�PH�EP���$Q���  �у�]� ��������U���SV��������؉]����   �} ��   �t��HH��p  j h�  V�҃��E��u
^��[��]� �MW3��}����������   �]��I �E�P�M�Q�MW������ta�u�;u�Y�I ������u�E�������L�;Ht-�t��Bl�S�@����QR�ЋD������t	�M�P�s���F;u�~��}��MG�}��>���;��v����]�_^��[��]� ^3�[��]� ��������������U����t�SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u�t��HH���  �'��u�t��HH���  ���ušt��HH���  S�ҋȃ��E��t�W�����t��HH���   h�  S3��҃����  ���_�u����    �t��Hl�U�B�IWP�ы�������   �t��F�J\�UP�A,R�Ѓ���t�K�Q�M�%����t��F�J\�UP�A,R�Ѓ���t�K�Q�M������E��;Pt&�F�t��Q\�J,P�EP�у���t	�MS������t��v�B\�M�P,VQ�҃���t�M�CP�����t��QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U��t��HH���   ]�������������̡t��PH���   Q��Y��������������U��t��HH���  ]��������������U��t���P���   V�uW�}���$V�����E������At���E������z����؋t��Q�B,���$V����_^]����������������U���0��t��U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١t��]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U��t��HH�]��U��t��H@�AV�u�R�Ѓ��    ^]�������������̡t��HH�h�  �҃�������������U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��HH�Vh  �ҋ�������   �EPh�  �`�������t]�t��QHj P���   V�ЋMQh(  �6�������t3�t��JH���   j PV�ҡt����   �B��j j���Ћ�^]át��H@�QV�҃�3�^]�������U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��HH�Vh�  �ҋ�����u^]át��HH�U�E��  RPV�у���u�t��B@�HV�у�3���^]�������U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��HH�I]�����������������U��t��H@�AV�u�R�Ѓ��    ^]��������������U��t��PH�EPQ���  �у�]� �U��t��PH�EPQ���  �у�]� ̡t��PH���  Q�Ѓ�������������U��t��HH���  ]��������������U��t��E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡t��PH���  Q�Ѓ�������������U��t��PH�EP�EPQ���  �у�]� ������������̡t��PH��  Q�Ѓ�������������U��t��PH�EP�EP�EPQ���  �у�]� ��������̡t��PH���  Q�Ѓ������������̡t��PH���  Q�Ѓ�������������U��t��PH�EPQ��  �у�]� �U��t��PH�EPQ��  �у�]� ̋������������������������������̡t��HH���  ��U��t��HH���  ]��������������U��t��PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U��t��PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡t��PH��,  Q�Ѓ�������������U��t��PH�EPQ��X  �у�]� ̡t��PH��\  Q�Ѓ�������������U��t��HH��0  ]��������������U��t���W���HH���   j h�  W�҃��} u�   _��]� Vh�  �������������   �t��HH���   j VW�҃��M������t��P�E�R0Ph�  �M����E�t��P�B,���$h�  �M��Ћt��Q@�J(j �E�PV�у��M�����^�   _��]� ^3�_��]� �����U��S�]�; VW��u7�t��U�HH���   RW�Ѓ���u�t��QH���   jW�Ѓ���t�   �����   �t��QH���   W�Ѓ��} u(�t��E�QH�M���  P�ESQ�MPQW�҃��B�u��t;�t��U�HH�ER�USP���  VRW�Ћt����   �B(�����Ћ���uŃ; u�t��QH���   W�Ѓ���t3���   �W��u1�t��QH���   �Ћt��E�QH���   PW�у�_^[]� �t��BH���   �у��} u0�t��M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� �t��QH�h  �Ћ؃���u_^[]� �t����   �u�Bx���Ћt����   P�B|���Ѕ�tU�t��E�QH�MP�Ej Q���  VPW�у���t�t����   �ȋBHS�Ћt����   �B(���Ћ���u�_^��[]� ��������������U��EV���u�t��HH���  �'��u�t��HH���  ���u�t��HH���  V�҃���u3�^]� P�EP���>���^]� ���������U���D�t��HH���   S�]VWh�  S�ҋ�t��HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��.
  �t����   �B���Ћt�=�  ��  �QH���   Wh:  S�Ћt��QH�E����   h�  S�Ћt��QHW�����   h�  S�uԉ}��Ћt��QH�E苂  S�Ћt��QH�EЋ��  S�Ѓ�(�E��E��}��~~�M���M�I �MЅ�tMj�W�qO  ���t@�@�Ẽ|� �4�~����%�������;�u/���Y  ;E�~�E؋��aY  E���E�;Pu�E���E��E�G;}�|��}� tv�u�j S�����������  ���������tV���q����}�;�uK�t��H���  �4�h�}��h�  V�҃��E���N  �M�PVP�}���P�'`  ����}ܡt��H���  �4�h�}��h�  V�҃��E����  �M�3�;�t;�tVQP�ت  ���E�;�~-�t��Qh�}��h�  P���   �Ѓ��E�;���  �t��E��QH��  j�PS�у�����  �u�;�tjS���������{  ��������E���}�t��BH���   Wh�  S�у�3�9}ԉE�}��`  �}���}Ȑ�MЅ��R  �U�j�R�zM  ����>  �M̍@�|� ���]�~����%�������9E���  ���mW  �E�3�3�9C�E܉M���   ��$    �����������tk�]��}������������ϋ9�<��}�@�҉��y�]��|��]�@@�z�<��y�]��|��]�@@�z�<��I�}��]�@���M��}�@����@�M�A;K�M��t����E؅��9  �+U�j��PR�M���9  �M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$��i�U����4�"�M����t��U����t�
�M����t�M���;]�|��E܃�F;]؉M��	����U�;U��
  �U�R��o���E�P��o���M�Q�o����_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���P�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@��;EԉE��}�������U�R�m���E�P�m�����  ���   �B����=  ��  �t��QH���   j h(  S�Ћt��QH�����   h(  S�ЋЃ�3��U؅�~'����    �ǅ�t�|� t�4N��tN�@;�|�u��u܋t��Q���  �4v�h�}��hK  V�Ѓ��E�����   �M��t��tVQP��  ���u؋t��Q���  �h�}��hP  V�Ѓ��E���tP��t��tVWP覤  ���M����+t��RH��PQ�E���   S�Ѓ���u�M�Q�bl���U�R�Yl����_^3�[��]át��HH���   j h�  S�҉E��t��HH���   j h(  S��3�3���3�9]؉E��}ĉ]��7  �U��څ��  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�F@F����;�|��}ă|� ts�U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�F�v�Ћ��A�B�A�B�A�B�A�B�I�J�U�F<ډ}�C;]؉]�������M�3�3�;�~�U����$    ��t���   @;�|��U�R�j�����E�P�j����_^�   [��]��c�c�cd������������U��E� �M+]� ���������������U��V��V��}�t��Hl�AR�Ѓ��Et	V�Tm������^]� ����������h��Ph�f �.  ���������������U���Vh��h�   h�f ���S.  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh��h�   h�f ����-  ����t���   ��t�M�UQ�MRQ����^]� U���Vh��h�   h�f ���-  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh��h�   h�f ����,  ����t���   ��t�M�UQ�MRQ����^]� U��Qh��h�   h�f �,  ����t���   �E���t�EP�U�����]��Pv��]�������������U���h��h�   h�f �f,  3Ƀ�;�tK9��   tC�E���   ���M��$Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]ËE�   � �  �P�P�H�H�H��]��U��h��h�   h�f ��+  ����t���   ��t]��]����U��h��h�   h�f �+  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h��h�   h�f �I+  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h��h�   h�f ��*  ����t���   ��t]��3�]��U���Vh��h�   h�f �*  ����tZ���   ��tP�M�UWQR�M�Q�Ћt��u���B�HV�ыt��B�HVW�ыt��B�P�M�Q�҃�_��^��]át��H�u�QV�҃���^��]����������h��h�   h�f �*  ����t���   ��t��3��������U��h��h�   h�f ��)  ����t���   ��t]��]����U��VWh��h�   h�f �)  ������tb���    tY�E �M�UP�t�Q�HR�Q����V�ҡt��H�A�UVR�Ћ��   ���ыt����B�P�MQ�҃� ��_^]át��H�A�UR�Ѓ�_3�^]���U��VWh��h�   h�f �)  ������tb���    tY�E �M�UP�t�Q�HR�Q����V�ҡt��H�A�UVR�Ћ��   ���ыt����B�P�MQ�҃� ��_^]át��H�A�UR�Ѓ�_3�^]���U���Vh��h�   h�f �u(  ����tZ���   ��tP�M�UWQR�M�Q�Ћt��u���B�HV�ыt��B�HVW�ыt��B�P�M�Q�҃�_��^��]át��H�u�QV�҃���^��]����������U���Vh��h�   h�f ��'  ����tS���   ��tI�MWQ�U�R�Ћu���t��H�QV�ҡt��H�QVW�ҡt��H�A�U�R�Ѓ�_��^��]Ët��Q�u�BV�Ѓ���^��]����������������U���Vh��h�   h�f �5'  ����tS���   ��tI�MWQ�U�R�Ћu���t��H�QV�ҡt��H�QVW�ҡt��H�A�U�R�Ѓ�_��^��]Ët��Q�u�BV�Ѓ���^��]����������������U��h��h�   h�f �&  ����t���   ��t]��]����U��h��h�   h�f �i&  ����t���   ��t]��]����U��M��U+u&�A+Bu�A+Bu�A+Bu�A+Bu�A+B]����������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���h���   h�   h�f �E��  �E��E��E�    �E�    �E�    ��#  ����t���   ��t	�M�Q�Ѓ��UR�E�P��������]��U��E��u����MP�EPQ裣����]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h~j;h��j��b������t
W�������3��F��u_^]� �~ t3�9_��^]� �t��H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   �t��H<�Q��3Ʌ����^��������������̃y t�   ËA��uËt��R<P��JP�у��������U����u�t��H�]� �t��J<�URP�A�Ѓ�]� ���������������U�졐���u�t��H�]Ët��J<�URP�A�Ѓ�]�U�졐���$V��u�t��H�1��t��J<�URP�A�Ѓ����t��Q�J�E�SP�ыt��B�P�M�QV�ҡt��H�A�U�R�Ћt��Q�Jj j��E�h\~P�ыt��B�@@�� j �M�Q�U�R�M��Ћt��Q�J���E�P���у���[t.�t��B�u�HV�ыt��B�P�M�Q�҃���^��]át��P�E��RHjP�M��ҡt��P�E�M��RLj�j�PQ�M��ҡt��H�u�QV�ҡt��H�A�U�VR�Ћt��Q�J�E�P�у���^��]���������������U�졐���$SV��u�t��H�1��t��J<�URP�A�Ѓ����t��Q�J�E�P�ыt��B�P�M�QV�ҡt��H�A�U�R�Ћt��Q�Jj j��E�h\~P�ыt��B�@@�� j �M�Q�U�R�M��Ћt��Q�J���E�P���у���t/�t��B�u�HV�ыt��B�P�M�Q�҃���^[��]át��P�E��RHjP�M��ҡt��P�E�M��RLj�j�PQ�M��ҡt��H�A�U�R�Ћt��Q�Jj j��E�h\~P�ыt��B�@@��j �M�Q�U�R�M��Ћt��Q�J���E�P���у����3����t��P�E��RHjP�M��ҡt��P�E�M��RLj�j�PQ�M��ҡt��H�u�QV�ҡt��H�A�U�VR�Ћt��Q�J�E�P�у���^[��]����������������U�졐���$SV��u�t��H�1��t��J<�URP�A�Ѓ����t��Q�J�E�P�ыt��B�P�M�QV�ҡt��H�A�U�R�Ћt��Q�Jj j��E�h\~P�ыt��B�@@�� j �M�Q�U�R�M��Ћt��Q�J���E�P���у���t/�t��B�u�HV�ыt��B�P�M�Q�҃���^[��]át��P�E��RHjP�M��ҡt��P�E�M��RLj�j�PQ�M��ҡt��H�A�U�R�Ћt��Q�Jj j��E�h\~P�ыt��B�@@��j �M�Q�U�R�M��Ћt��Q�J���E�P���у����3����t��P�E��RHjP�M��ҡt��P�E�M��RLj�j�PQ�M��ҡt��H�A�U�R�Ћt��Q�Jj j��E�h\~P�ыt��B�@@��j �M�Q�U�R�M��Ћt��Q�J���E�P���у���������t��P�E��RHjP�M��ҡt��P�E�M��RLj�j�PQ�M��ҋu�E�P��裓���t��Q�J�E�P�у���^[��]�������U�졐���$SV��u�t��H�1��t��J<�URP�A�Ѓ����t��Q�J�E�P�ыt��B�P�M�QV�ҡt��H�A�U�R�Ћt��Q�Jj j��E�h\~P�ыt��B�@@�� j �M�Q�U�R�M��Ћt��Q�J���E�P���у���t/�t��B�u�HV�ыt��B�P�M�Q�҃���^[��]át��P�E��RHjP�M��ҡt��P�E�M��RLj�j�PQ�M��ҡt��H�A�U�R�Ћt��Q�Jj j��E�h\~P�ыt��B�@@��j �M�Q�U�R�M��Ћt��Q�J���E�P���у����3����t��P�E��RHjP�M��ҡt��P�E�M��RLj�j�PQ�M��ҡt��H�A�U�R�Ћt��Q�Jj j��E�h\~P�ыt��B�@@��j �M�Q�U�R�M��Ћt��Q�J���E�P���у���������t��P�E��RHjP�M��ҡt��P�E�M��RLj�j�PQ�M���j h\~�M��B����t��P�R@j �E�P�M�Q�M��҅��t��H�A�U�R���Ѓ���t/�t��Q�u�BV�Ћt��Q�J�E�P�у���^[��]Ët��M��B�PHjQ�M��ҡt��P�E�M��RLj�j�PQ�M��ҋu�E�P���k����t��Q�J�E�P�у���^[��]���������������U��t��H<�A]����������������̡t��H<�Q�����V��~ u>���t�t��Q<P�B�Ѓ��    W�~��t���
���W�$W�����F    _^��������U���V�E�P���>�����P��������M���������^��]��̃=�� uK�����t�t��Q<P�B�Ѓ����    �����tV������V�V�������    ^������������U���8�t��H�AS�U�V3�R�]��Ћt��Q�JSj��E�h`~P�ыt��B<�P�M�Q�ҋ�t��H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��  �M�Q�U�R�M���  ����   W�}�}���   �t����   �U��ATR�Ћ�����tB�t��Q�J�E�P���у��U�Rj�E�P��輎���t��Q�ȋBxW���E���t�E� ��t�t��Q�J�E�P����у���t�t��B�P�M�Q����҃��}� u"�E�P�M�Q�M��/  ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3ۉ]�;�u_�t��H�A�U�R�Ћt��Q�JSj��E�h`~P�ыt��B<�P�M�Q�ҋ�t��H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��!  �M�Q�U�R�M��q  ���p  W�}��I �E����   �t����   �U��ATR�Ћ�������   �t��Q�J�E�P���ыt��B���   ���M�Qj�U�R���Ћt��Q�J���E�P�ыt��B�P�M�QV�ҡt��H�A�U�R�Ћt��Q�Bx��W�M����E��t�E ��t�t��Q�J�E�P����у���t�t��B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*�t����   P�BH�Ћt��Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��s  �EP�M�Q�M�u��u�  ����   �u���E���tA��t<��uZ�t����   �M�PHQ�ҋt��Q���ȋBxV�Ѕ�u-�   ^��]Ët����   �E�JTP��VP�[�������uӍUR�E�P�M��4  ��u�3�^��]����������V��~ u>���t�t��Q<P�B�Ѓ��    W�~��t�������W��Q�����F    _^�������̋�� p~���������p~���������̅�t��j�����̡t��P��  ��t��P��(  ��U��t��P��   ��V�E�P�ҋuP��������M��2�����^��]� ��������̡t��P��$  ��U��t��H��  ]��������������U��t��H���  ]�������������̡t��H��  ��U��t��H���  ]��������������U��t��H��x  ]��������������U��t��H��|  ]�������������̡t��H��d  ��U��t��H��p  ]��������������U��t��H��t  ]��������������U���EV���p~t	V�P������^]� �������������̸   � �������̸   @� �������̸   � �������̸   � ��������U��t��H�QV�uV�҃���^]� �3�� �����������3�� �����������3�� �����������U����   h�   ��@���j P�Td  �M�Eh�   ��@���R�M��MPQjǅ`���    �yx���� ��]���U����   V�u��u3�^��]�h�   ��@���j P��c  �M�U�Eh�   �M���@���Q�U��U��@����ERPj��`���ǅD������E�P��E����E����E� ��E�Ў�E�`��E����E�����w���� ^��]������U���   SV�u(3ۉ]���u�t��H�A�UR�Ѓ�^3�[��]Ët��Q�B<W�M3��Ѕ��'  �8  �E���tq�MQ�M��i���Wht~�M��ۆ��P�M��R����u�Wj��U�R�E�P��\���Q�_?������P��x���R������P�E�P�������P����9  �E���t�E� �� t�M�����p�����t��x�������]�����t��\�������J�����t�M̃���:�����t�t��Q�J�E�P����у���t�M������}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R�7  ����E$�M�UVP�Ej QRP����������t��Q�J�EP�у���_^[��]���������������̋�`����������̋�`����������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V����5  �����   �ESP�M��Ⱦ���t��Q�J�E�P�ыt��B�Pj j��M�ht~Q�҃��E�P�M�茾��j j��M�Q�U�R��d���P�T�����P�M�Q�G�����P�U�R�:������P�7  ���M���������M�蹾����d���设���M�覾���t��H�A�U�R�Ѓ��M�芾����[t	V�/5  ����^��]� ���U��EVP����?  �����^]� �����Q��4  Y���������U��E�M�U�H4�M�P �U��M�@���@8P��@<���@@���@D���@H���@L`��@P ��@lp��@X���@\0��@`���@d���@TЎ�@h���@p��@t@��P0�H(�@,    ]��������������U���   h�   ��`���j P�^  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�r����8��]��������������̋�`<����������̋�` ����������̋�`0����������̋�`@����������̋�`����������̋�`����������̋�`$����������̋�`4����������̋�`����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U��E��u�E�M�������   ]� �����������U��EHV����   �$�(��   ^]á��@�����uT�EP觺����=�.  }�����^]Ëu��t�hx~jmh��j�H������t ��譺�������tV��輾���   ^]����    �   ^]ËM�UQR�Ÿ���������H^]�^]�p����-��u.蒸���}��������t���,���V�FG�������    �   ^]Ã��^]ÍI @�ُ��8����U���EV���V��������Au�t��H��0  h�~j,�����^��^]� �����U���W������G���U���}������A�  ������A��   � ������AuR������AuKV���[y  ���Ty  �ȅ�u��^����__��]Ëƙ����ʅ�u�u��E�^������__��]���������Au������=��������Au6�����������U������G�����_��������Au�����U����_�
����������]  �E����U����������A{���������__��]�������������__��]����U���0V�E��������At���(������Au������|����$��v  ����|���^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3����;���W���$���v  ��E����$�lv  �V����������Au�t��H��0  h�~j�����^����_u������������^]� ���U������EV�ы�������z!�t��؋H��0  h�~j5�����U������$��u  �]��F�$��u  �}��$��u  ��E�$�u  �^�����&���^��]� ���������������U��t����   �BXQ�Ѓ���u]� �t��Q|�M�RQ�MQP�҃�]� ���U��t����   �BXQ�Ѓ���u]� �t��Q|�M�R8Q�MQP�҃�]� ���U��EV��j ��t��Qj j P�B�ЉF����^]� ��̡t�Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� �t��Q�MP�EP�Q�JP�у��F�   ^]� ����U��M��P]����U��M��P]����U��M��P]����V���<�F    �t��HP�h��Vh��h���҉F����^����������̃y �<u�t��PP�A�JP��Y��U��A��u]� �t��QP�M�Rj Q�MQP�҃�]� ��U��A��t�t��QP�M�RQP�҃�]� ������������U��A��t�t��QP�M�RQP�҃�]� �����������̡t��HP���   ��U��t��HP���   ]�������������̡t��HP�QP�����U��t��HP�AT]����������������̋��     �@    �V����t)�t��QPP�BL�Ћt��QP��J<P�у��    ^�������������U��SV�ً3�W;�t�t��QPP�B<�Ѓ��3�s�}�Eh��W�C�t��QP�J8h��h��P�EP�у�9u�~M�I ���z u!���@   �t��QP���H�RQ�҃��t��HP��A@VR�Ћ�F��;u�A|�3�9_^��[]� ��������U��SVW��3�9w~<�]�t��HP��A@VR�Ѓ���t-�t��QPj SjP�B�Ѓ���tF;w|�_^�   []� �t��QP��JLP�у�_^3�[]� �����������̡t��PP��JDP�у�������������̡t��PP��JHP��Y��������������̡t��PP��JLP��Y���������������U��U�E�@R�URP�I���]� �����U��V��~ �<u�t��HP�V�AR�Ѓ��Et	V��>������^]� ����U��E�M�UP��P�EjP��l����]��������������̸   �����������U��V�u��t���u6�EjP��l������u3�^]Ë���m����t���t��U3�;P��I#�^]�������U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �������������U��V�u�F��F�����������������|q  ����������D�Ez��^��P�X]��������������N�X�N^�X]��������P�P�P�P �P(�P0�P8�P@�PH�PP�PX����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��5�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A �A�A(�A�����������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E������X�X]� ̋�3ɉ�H�H�H�V��V�0���FP�0��3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  S�]���q  ��؋�U��M�U�>�U��@�����@�U��@�B�@�������@���@�   ;����U��p  �w�����  �w�������F�B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]؋�R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ɍU��R�[�[������E��KH��P�E�SL��H�щKP�P�ST�H�KX�P�����S\��z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����M��}������3�3����u��u�|+�A�����B�4�u�0u��u�p�����u�u�U�E;�}�Q���E����U��U��1���@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���@�D��KX�@�U�����]��C���@�K0���@�KH���C ��C�@�K8���@�KP���C(��C�C@�H���@3����KX���U��r  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�E�KX@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������]��E�E����]���E����]��E׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���@�KX���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���@�   �KXE)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� ������������h��Ph_� �������������������h��jh_� ��������uË@����U��V�u�> t/h��jh_� �c�������t��U�M�@R�Ѓ��    ^]���U��Vh��jh_� ���)�������t�@��t�MQ����^]� 3�^]� �������U��Vh��jh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh��jh_� ����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��jh_� ���Y�������t�@��t�MQ����^]� 3�^]� �������U��Vh��j h_� ����������t�@ ��t�MQ����^]� 3�^]� �������U��Vh��j$h_� �����������t�@$��t�MQ����^]� 2�^]� �������Vh��j(h_� ����������t�@(��t��^��3�^������Vh��j,h_� ���l�������t�@,��t��^��3�^������U��Vh��j0h_� ���9�������t�@0��t�MQ����^]� 3�^]� �������U��Vh��j4h_� �����������t�@4��t�M�UQR����^]� ���^]� ��Vh��j8h_� ����������t�@8��t��^��3�^������U��Vh��j<h_� ����������t�@<��t�MQ����^]� ��������������U��Vh��j@h_� ���I�������t�@@��t�MQ����^]� ��������������U��Vh��jDh_� ���	�������t�@D��t�MQ����^]� 3�^]� �������U��Vh��jHh_� �����������t�@H��t�MQ����^]� ��������������Vh��jLh_� ����������t�@L��t��^��3�^������Vh��jPh_� ���\�������t�@P��t��^��3�^������Vh��jTh_� ���,�������t�@T��t��^��^��������Vh��jXh_� �����������t�@X��t��^��^��������Vh��j\h_� �����������t�@\��t��^��^��������U��Vh��j`h_� ����������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh��jdh_� ���Y�������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh��jhh_� ����������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh��jlh_� �����������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��jph_� ���y�������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh��jth_� ���9�������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh��jxh_� �����������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh��j|h_� ����������t�@|��t�MQ����^]� 3�^]� �������U��Vh��h�   h_� ���v�������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h_� ���&�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh��h�   h_� �����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh��h�   h_� ���f�������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h�   h_� ����������t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   h_� �����������t���   ��t�MQ����^]� ��������U��Vh��h�   h_� ����������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h_� ���F�������t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E����������m������U�_��^�U�[���U������������������������6Y  ����������D�Ez����P�X��]� �������E�����E����X�M��X��]� �����U���@� |�A���E�    �����]��]��]���{�������]��]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P�q����F�@��R�M��_����~���Q�M��M����v;�t�v��P�M��7����M����m��M�u�_^[�M�UQR�M��������]� ��������������̋Q3���|�	��t��~�    t@����u��3���������U��QV�u;��}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��|+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~#V�1�d$ ���   @u	�����t@����u�^���̋QV3���~�	�d$ ����ШtF����u��^���������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%���;��E���}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$�H��E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� �������3�����U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V����FP���3����F�F^��U��SV��WV�����^S�����E3����~�~;�t_�t��Q���   hP��jIP�у��;�t9�}��t;�t��B���   hP��    jNQ�҃����uV�{����_^3�[]� �E�~_�F^�   []� ����������U��SV��WV�B���^S�9���}3Ƀ��N�N;���   9��   �G;���   �t��Q���  hP��jlP�у����t=� t@�G��t9�t��JhP��    ���  jqR�Ѓ����u������_^3�[]� �O�N�G�Q��    R�F�QP�  �����t�N�WP��QPR�x  ��_^�   []� ���������U��SV��WV�B���~W�9��3Ƀ��N�N9M��   �E;���   ��    �t��H���  hPh�   S�҃����t=�} tH�E��tA�t��Q���  hP��h�   P�у����u������_^3�[]� �U�V�,�F   �t��H���  hPh�   j�҃����t��E�M�F�PSPQ�q  �E����t!�V�?�W�RWP�U  ��_^�   []� ��M�_^�   []� ���U��Q�A�E� ��~LS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U�����u�_^[�E��Ћ�]� ���������U��S�]V��3�W�~���F�F�CV;C��   ���W�~��3��F�F�t��Q���   hPjIj�Ѓ������   �t��Q���   hPjNj�Ѓ����uV�&����_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� ����W����3��F�F�t��B���   hPjIj�у����t[�t��B���   hPjNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP��������^]� ����������U��U��t�M��t�E��tPRQ��J  ��]�����������̡t��H���   ��U��t��H���   V�u�R�Ѓ��    ^]����������̡t��P���   Q�Ѓ�������������U��t��P�EPQ���   �у�]� ̡t��H�������U��t��H�AV�u�R�Ѓ��    ^]��������������U��t��H�AV�u�R�Ѓ��    ^]��������������U��t��P��Vh�  Q���   �E�P�ыt����   �Q8P�ҋ�t����   ��U�R�Ѓ���^��]��������������̡t��P�BQ�Ѓ����������������U��t��P�EPQ�J\�у�]� ����U��t��P�EP�EP�EP�EP�EPQ���   �у�]� �U��t��P�EP�EP�EP�EPQ�JX�у�]� �������̡t��P�B Q��Y�U��t��P�EP�EP�EP�EPQ���   �у�]� �����U��t��P�EP�EP�EPQ�J�у�]� ������������U��t��H��   ]��������������U��t��P�R$]�����������������U��t��P��x  ]�������������̡t��P��|  ��U��t��P�EP�EP�EP�EPQ�J(�у�]� ��������U��t��P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U��t��P�EP�EP�EP�EPQ�J,�у�]� ��������U��t�V��H�QWV�ҋ��t��H�QV�ҋt��Q�M�R4Q�MQ�MQOWHPj j V�҃�(_^]� ���������������U��t��P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U��t��P�EP�EPQ�J@�у�]� U��t��P�EPQ�JD�у�]� ���̡t��P�BLQ�Ѓ���������������̡t��P�BLQ�Ѓ���������������̡t��P�BPQ�Ѓ����������������U��t��P�EPQ�JT�у�]� ����U��t��P�EPQ�JT�у�]� ����U��t��P�EP�EPQ���   �у�]� �������������U��t��P�E���   ��VP�EPQ�M�Q�ҋu�    �F    �t����   j P�BV�Ћt����   �
�E�P�у� ��^��]� ������̡t��P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡t��H�������U��t��H�AV�u�R�Ѓ��    ^]��������������U��t��P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U��t��P�EPQ�J�у�]� ���̡t��P�BQ��Y�U��t��P�EP�EPQ�J�у�]� U��VW���t����M�U�x@�EPQR���^����H ���_^]� �U��VW���D����M�U�xD�EPQR���.����H ���_^]� �V�������xH u3�^�W�������΍xH������H �_^�����U��V�������xL u3�^]� W���м���M�U�xL�EPQR��躼���H ���_^]� �������������U��V��蕼���xP u���^]� W�������M�U�xP�EP�EQRP���e����H ���_^]� ��������U��V���E����xT u���^]� W���/����M�xT�EPQ�������H ���_^]� U��V�������xX u���^]� W�������xX�EP�������H ���_^]� ����U���S�]VW���t.�M�趢����读���xL�E�P��衻���H ��ҍM������}��tZ�t��H�A�U�R�Ћt��Q�J�E�WP�ыt��B�P�M�Q�҃����I����@@��t�t��QWP�B�Ѓ�_^[��]� ������U��V�������x` u
� }  ^]� W��������x`�EP�������H ���_^]� ��U��VW���Ժ���xH�EP���ƺ���H ���_^]� ���������U��SVW��裺���x` u� }  �#��菺���x`�E���P���|����H ��ҋ��t��H�]�QS�҃�;�A�t��H�QS�҃�;�,���?����M�U�xD�EPQSR���(����H ���_^[]� _^�����[]� ��������������U��V��������xP u
�����^]� W���ݹ���M�U�xP�EP�EQ�MR�UPQR��軹���H ���_^]� ��������������U��V��蕹���xT u
�����^]� W���}����M�xT�EPQ���k����H ���_^]� ��������������U��V���E����xX tW���7����xX�EP���)����H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u���  ����t.�E�;�t'�t��J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡t��H��   ��U��t��H��$  V�u�R�Ѓ��    ^]�����������U��t��UV��H��(  VR�Ѓ���^]� �����������U��t��P�EQ��,  P�у�]� �U��t��P�EQ��,  P�у����@]� �����������̡t��H��0  ��t��H��4  ��t��H��p  ��t��H��t  ��U��E��t�@�3��t��RP��8  Q�Ѓ�]� �����U��t��P�EPQ��<  �у�]� �U��t��P�EP�EP�EPQ��@  �у�]� ���������U��t��P�EP�EPQ��D  �у�]� �������������U��t��P�EPQ��H  �у�]� �U��t��P�E��L  ��VWPQ�M�Q�ҋu���t��H�QV�ҡt��H�QVW�ҡt��H�A�U�R�Ѓ�_��^��]� ��������������̡t��P��T  Q�Ѓ�������������U��t��P�EPQ��l  �у�]� ̡t��P��P  Q�Ѓ�������������U��t��P�EPQ��X  �у�]� ̡t��H��\  ��U��t��H��`  V�u�R�Ѓ��    ^]�����������U��t��P�EP�EP�EP�EP�EPQ��d  �у�]� �U��t��P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w����y����3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7��迴���xP t$S��豴��j j �XPj�FP��蝴���H ���[�    �~` t�t��H�V`�AR�Ѓ��F`    _^������������U��SV��Fx�t��Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR�3������u#���h��t��H��0  h  �҃��E�~P���||���j j jW�����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    �t��Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ��i����F|��u�E�~x��t�    �F`_^]� �M�Fx������t�3�_^]� U��QVW�}����>  �t��H�QhV�҃����t�u"�H��0  h�h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���  �EF;u�|�UR� ����_�   ^��]� �������������U��QVW�}����~  �t��H�QhV�҃����t�u"�H��0  h�h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'���t��QP�Bh�Ѓ���t�M��R���,  F;u�|ʍEP������_�   ^��]� �������������h�h�   h��h�   �w������t�������3��������V���(����N^�ov�����������������U��VW�}�7��t��������N�Cv��V�]�����    _^]�h��Ph�f �������������������U��h��jh�f �l�������t
�@��t]�����]�������U��Vh��jh�f �;���������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�Zu���E�NP�у�4�M���u����^]ÍM�wu�����^]��U��h��jh�f ���������t
�@��t]��3�]��������U��h��jh�f ��������t�x t�P]��3�]������V��FW��u�~��N�<��u�< ��u_3�^át��H�F��  h�j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� }(�V;Vu��������t�F�N��    �F9~|؋V;Vu���������t��F�N�U���F_�   ^]� ��������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T����H;ǉ�F�M���F_�   ^]� ����U��E��|2�Q;�}+J;Q}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�����3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�L������3����_�F�F^��������������U���SV�uW���^S�}�����3���F�F�O�N�W���V9G�E~|��I �O���F�U�9FuL��u�~��~��t���< ��tY�t��H���  h�j8��    RP�у���t0�~�}���V��M����E�F@;G�E|�_^�   [��]� _^3�[��]� U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|���P�����_^]� �U����E�Qj�E��ARP�M��E�T��������]� �����U����Q�Ej�E��A�MRPQ�M��E�T�������]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q����t!�A��t�B�A�Q�P�A    �A    �̋�� \��@��HV3��q�q�P�r�r���p�p�p�P�H^������V���\������F3��F�;�t�N;�t�H�F�N�H�V�V�F�F�;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3���;�t�F;�t�A�F�N�H�V�V�Et	V��������^]� ������������U��V��W�~W�L��*���3����E��F�Ft	V�Q�����_��^]� ������U��V��������Et	V�)�������^]� ��U���V�u��u��=  �@�E��=  ���E�F�}� �E�u�E�H�����   �� ��   S�]W�   ;�s��uS�7  Y��u�   �F�Xt}��u�]��}���6  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPW�u�j �S6  ��$��u������E�t	�M����_[^�Ë�U��V��<  �@�u��<  jh   �F�-=  YY�F��th   �<6  P�v�,  ���F   ��"6  �f �F��^]Ë�Wh�����p��uV���V��  ���� �Y|�^��_�h���p��}V���V�  ���� �Y|�^Ë�U��E��V��}k���P�  Y��^]� ���}k���P�  YË�U���u�h0  Y��t]�=  ]ËI�w�����t�j���Ë�U��V��������EtV�����Y��^]� ��U��E���t�6�����t�j���]Ë�U��Qj �M��@���h(�������%(� Y�M��N����á(�Ë�U��=L� uh���L���  Y�E�(�]�j�-h�3>  j �M�������}�e� �w��GN���8 t�藷����t�j�����w��w�b  �M��Y�M�������I>  Ë�U��Qj �M�������ȋ j�$�������$���u�M������Ë�U��=$� uhd�����Yj����Y��t�$���M�H�3��$�]Ë�U��E�xP v�xTr�@@���@Pj �L  YY]�j�Ph�8=  ��u��F   3��E��F�F�F�Ehh��N�d��F�r9�����g=  � j�~h��<  ��u��d�V�E�   ����Yj j�N�!����v�(=  Ë�U��V�������EtV����Y��^]� j��h�<  �(�����u{P�M��2����(�!u�����uXj4�u���Y�ȉM��E���t
V�������3�V�E� ������N�F?   �$l��[1���Ή5,��~����,��D��M���M���������m<  Ë�U��E�xVWr�p��pj j �J  YY��u��r�}P�O<��0����tVj �~J  YY��u�h�P�OX��0��_^]Ë�U��VW���w ��vW�u�V�6����u�_^]� ��U��V�uWj ��������F��t�8P�k���Y�ǅ�u�F �f ��t�8P�Q���Y�ǅ�u�f  _^]Ë�U��V�u�~ v�F�����F���� V����Y�N$��tj�y��^]Ë�Vj�������P��2  YY��^Ë�V���6�0  �6�����YY^��1�.  Y��1�5  YË�U���V�u��u�7  �@�E��T7  ���E�F�}� �E�u�E�H�����   �� ��   S�]��   s!��uS��1  Y��u�   �F�X��   ��u�]��}��0  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPh   �u�j ��/  ��$��u������E�t	�M����[^�Ë�U��V�u���4���x���^]� �x��i4����U��V���x��V4���EtV�j���Y��^]� jD��h�I9  h���M��5���e� �E�P�M���3��hH��E�P�B  �jD��h�9  h���M��q5���e� �E�P�M��P���hл�E�P�
  ̋�U��V�u���B<���x���^]� ��U��USVW�ڋ�����   ��@t����t��3Ɂ�;���3�A;�t����@��u��������� u3��^��t%��t �uh���u�H  ����t	P�  Y���u��H�V�u�gH  ������t���tjj V�8  ����tV�ŋ�_^[]Ë�U���  ��3ŉE��Eh  Ph  ������Pj �K  ����t3���u�������uP��������M�3��  �Ë�U���u� p]Ë�U���u�$p]Ë�U���u�(p]Ë�U���u�,p]Ë�U�졌���u]�'6  �MH�������]������@�����t���������
r������̋L$WSV��|$��to�q��tU���L$���:�t��t���:�t
��u�^[_3�Ê��:�u�~��a��t(���:�u��A��t�f���:�t��3�^[_���J  �G�^[_Ë�^[_Ë�Q�<��*K  YË�U��V��������EtV����Y��^]� ��U��E��	Q��	P�dK  ��Y�Y@]� ��U��E��t���8��  uP�  Y]Ë�U��EV���F ��uc�SU  �F�Hl��Hh�N�;��t����Hpu�>9  ��F;��t�F����Hpu�M  �F�F�@pu�Hp�F�
���@�F��^]� ��U�����3ŉE�S3�V;�u�hX  j^SSSSS�0�e  ���5  �uW��W  YY;Er��ЋU��H;�u ��8t�<a|<z, �A8u�3���   j�p�   SSj�WVQR�D+  �ȃ�$�M�;�u��W  � *   ��W  � �   9Ms���W  j"�^���;�~Ej�3�X���r9�A=   w��W  ��;�t� ��  �P�   Y;�t	� ��  ���M�E���]�9]�u�nW  �    냋U�j�pQ�u�j�WV�pR�*  ��$��t�u��uW��   ������,W  j*Y����u������Y�ƍe�^[�M�3��  �Ë�U���W�u�M�������}�E�P�u�_����}� YY_t�M��ap��Ë�U��j �u�u������]Ë�U��S3�9�uA�E;�u�V  SSSSS�    �	  ��3��/��8t)�
��a|
��z�� �
B8u��Sj��u�X����E��[]Ë�U��MS3�VW;�t�};�w�;V  j^�0SSSSS�8	  �����0�u;�u��ڋъ�BF:�tOu�;�u�� V  j"Y�����3�_^[]�;�u���XV  �����������̋T$�L$��ti3��D$��u��   r�= t�}W  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�ø�O�P��T��F�X��F�\��F�`�<F�d��h�wO�l�XF�p��E�t�GEË�U�������rc  �} ���t��b  ��]���U��WV�u�M�}�����;�v;���  ��   r�= tWV����;�^_u^_]��c  ��   u������r*��$�����Ǻ   ��r����$����$�����$�X�����8�#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I ��������������x��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�`������$���I �Ǻ   ��r��+��$�d��$�`��t������F#шG��������r�����$�`��I �F#шG�F���G������r�����$�`���F#шG�F�G�F���G�������V�������$�`��I ��$�,�4�<�D�W��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�`���p�x������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ���` �` � P�Ë�U��S�]VW���P����t&P�\,  ��FV��  YY�G��t�3VP��������g �G   ��_^[]� ��U��S�]V���P��C�F���CWt1��t'P��+  ��GW�  YY�F��t�sWP�/������	�f ��F_��^[]� �y �P�t	�q��  YËA��u�X�Ë�U��V�EP�������p���^]� ��U��V�u���R����p���^]� �p�������U��V�������EtV����Y��^]� ��U��V���p��c����EtV�����Y��^]� ��U��V�uW3�;�u3��e9}u�O  j^�0WWWWW�  �����E9}t9urV�u�u�p  �����uW�u������9}t�9us�RO  j"Y����jX_^]�������������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[Ë�U��EVW3�;�tG9}u�nN  j^�0WWWWW�k  �����)9}t�9Es�IN  j"Y�����P�u�u�_�����3�_^]Ë�U��E���]Ë�U���(  ��3ŉE������� SjL������j P������������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������@pj ���<p��(���P�8p��u��uj�.]  Yh ��4pP�0p�M�3�[�����Ë�U���5����F  Y��t]��j��\  Y]����3�PPPPP�������Ë�U��� �EVWjY�x��}��E��E_�E�^��t� t�E� @��E�P�u��u��u��Dp�� jh��i  �u��tu�=�
uCj�^  Y�e� V�^  Y�E��t	VP��^  YY�E������   �}� u7�u�
j�}]  Y�Vj �5���Lp��u��K  ���HpP�K  �Y�ei  Ë�U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$����U��QQSVWd�5    �u��E���j �u�u��u�o �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�+v  �� �E�_^[�E���]Ë�U��V��u�N3�����j V�v�vj �u�v�u��u  �� ^]Ë�U���8S�}#  u����M�3�@�   �e� �E�����M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E��F  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M�����E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u�t  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����-���u�u  �M�N��k���M9H};H~���u	�M�]�u�} }ʋEF�0�E�;_w;�v�<u  ��k�E�_^[�Ë�U��EV�u��ME  ���   �F�?E  ���   ��^]Ë�U���*E  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V�E  �u;��   u��D  �N���   ^]���D  ���   �	�H;�t���x u�^]�t  �N�H�ҋ�U������e� �M�3��M�E��E�E�E@�E���M��E�d�    �E�E�d�    �uQ�u�t  �ȋE�d�    ����jh0��-e  3��}�3��u;���;�u ��G  �    WWWWW�����������   V�Wu  Y�}��F@uwV��y  Y���t���t�����ȃ��������P��A$u)���t���t�������������P��@$�t�OG  �    WWWWW�K������M��9}�u�Nx
��A��V�u  Y�E��E������   �E��d  ËuV�u  Y�jhP��)d  3��}�3��u;���;�u ��F  �    WWWWW�����������   V�St  Y�}��F@uwV��x  Y���t���t�����ȃ��������P��A$u)���t���t�������������P��@$�t�KF  �    WWWWW�G������M��9}�u!�Nx��E�����V�u�x  YY�E��E������   �E��zc  ËuV�t  YË�U��V�u�F@WuyV�!x  Y�P����t���t�ȃ��������������A$u&���t���t�ȃ������������@$�t�E  3�WWWWW�    �y���������JS�]���t=�F�u��y2�u.3�9~uV�y  Y�;Fu9~u@���F@�t8t@����[_^]È�F�F�����F��%�   ��jhp��,b  3�3�9u��;�u��D  �    VVVVV�����������+�u�\r  Y�u��u�u�����YY�E��E������	   �E��b  ��u�r  YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�v  YP�  ��;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�7v  P��  Y��Y��3�^]�jh���
a  3��}�}�j�V  Y�}�3��u�;5�
��   �����98t^� �@�tVPV�oq  YY3�B�U�������H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u����4�V�xq  YY��E������   �}�E�t�E��`  �j�kT  Y�jh���0`  3�9uu	V����Y�'�u�{p  Y�u��u����Y�E��E������	   �E��9`  ��u��p  Y�j�����Y�jhؼ��_  3ۉ]�3��u;���;�u �B  �    SSSSS�}���������   �E��t	;�t��@u�;�t��@u�}�G�=���v뷋}����uV��o  Y�]�V����V�6  YY�f�����N�Et���Fj_�-�E;�u W�  Y;�u����M����N  �	��   �N�~�F��^�E������	   �E��2_  ��u�o  YË�U���SVW3�9}t$9}t�u;�u�A  WWWWW�    ������3�_^[�ËM;�tڃ��3��u9Ew͋}�}�F  �M��}��t�F�E���E�   ����   �N��  t/�F��t(��   ��;�r��W�u��6��
  )~>��+�}��O;]�rO��tV�S���Y��u}�}� ��t	3ҋ��u�+�W�u�V�s  YP�|  �����ta��;�w��M�+�;�rP�}��)�E�� VP�s  YY���t)�E��FK�E����E�   ���A����E������N ��+�3��u������N �E���jh���t]  3�9ut)9ut$3�9u��;�u �@  �    VVVVV������3��]  ��u�m  Y�u��u�u�u�u�=������E��E������   �E����u��m  YË�U��W3�9}u�?  WWWWW�    ����������AV�u;�u�?  WWWWW�    �����������u��  Y�ȉ#ʃ���V;�t3�^_]Ë�U��V�u�F��u�@?  �    ����g���}�FuV�S�  E�e YV�����FY��y����F��t�t�   u�F   �u�uV�,q  YP�0�  3Ƀ������I��^]�jh���[  3�3�9u��;�u�>  �    VVVVV����������>�};�t
��t��u��u�l  Y�u�W�u�u�������E��E������	   �E���[  ��u�Yl  YË�U��V3�9uu�4>  VVVVV�    �0����������E;�t�V�p�0�u�p�  ��^]Ë�U��SV�uW3����;�u��=  WWWWW�    ���������B�F�t7V�:���V����z  V� p  P��  ����}�����F;�t
P�&���Y�~�~��_^[]�jh8��Z  �M��3��u3�;���;�u�e=  �    WWWWW�a����������F@t�~�E��Z  �V��j  Y�}�V�*���Y�E��E������   �ՋuV�!k  YË�U��Q�e� S�]��u3��   W��ru�{���vn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9}�r��?�@��I��F�@��I��<�@��I��2�@��I��(�M�E����t:u@A�E�9]�r�3�_[��� �	+����U���u�Tp��u�Hp�3���tP�N<  Y���]�3�]Ë�U��� WV�j  3�Y;�u�<  WWWWW�    �����������49}t޹����E�I   �u�u��M�;�w�E��u�E��u�uP�U��_�Ë�U��V�u�EPj �uh��z�����^]Ë�U��j
j �u�X�  ��]Ë�U��EVW��u|P�K  Y��u3��  �j9  ��u�K  ���ś  �\p��~�  �����j  ��}��5  ��詙  ��| �(�  ��|j ���  Y��u����   ��l  ��3�;�u19=��~����9=�u舖  9}u{��l  �5  �K  �j��uY�<5  h  j�  ��YY;��6���V�5���5T��4  Y�Ѕ�tWV�u5  YY�Xp�N���V�����Y�������uW��7  Y3�@_^]� jhX��vW  ����]3�@�E��u9����   �e� ;�t��u.�����tWVS�ЉE�}� ��   WVS�r����E����   WVS覆���E��u$��u WPS蒆��Wj S�B��������tWj S�Ѕ�t��u&WVS�"�����u!E�}� t�����tWVS�ЉE��E������E���E��	PQ葛  YYËe��E�����3���V  Ë�U��}u茛  �u�M�U�����Y]� ��������̃=�� ���  ���\$�D$%�  =�  u�<$f�$f��f���d$���  � �~D$f(��f(�f(�fs�4f~�fT��f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�L�  ���D$��~D$f��f(�f��=�  |!=2  �fT���\�f�L$�D$����f�ЁfVЁfT��f�\$�D$���������������̃= t-U�������$�,$�Ã= t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$��jhx��yT  �e� �u;5�
w"j�jI  Y�e� V�qQ  Y�E��E������	   �E��T  �j�eH  YË�U��V�u�����   SW�=`p�=�� u���  j�F�  h�   �H�  YY��
��u��t���3�@P���uV�S���Y��u��uF�����Vj �5���׋؅�u.j^9@�t�u�֞  Y��t�u�{����W6  �0�P6  �0_��[�V诞  Y�<6  �    3�^]��5L��70  Y��t��j蒜  jj �  ����  ��U��WV�u�M�}�����;�v;���  ��   r�= tWV����;�^_u^_]��D  ��   u������r*��$����Ǻ   ��r����$���$����$�(���#ъ��F�G�F���G������r���$���I #ъ��F���G������r���$���#ъ���������r���$���I �xph`XPH�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�0�����$���I �Ǻ   ��r��+��$�4�$�0�Dh��F#шG��������r�����$�0�I �F#шG�F���G������r�����$�0��F#шG�F�G�F���G�������V�������$�0�I ����'�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�0��@HXl�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U��QSVW�5���,  �5�����}��,  ��YY;���   ��+ߍC��rwW�Q�  ���CY;�sH�   ;�s���;�rP�u���  YY��u�G;�r@P�u���  YY��t1��P�4��+  Y����u�+  ���V�+  Y����EY�3�_^[�Ë�Vjj �G  ��V�h+  ����������ujX^Ã& 3�^�jh����N  �B�  �e� �u�����Y�E��E������	   �E�� O  ��!�  Ë�U���u���������YH]�������������̺@��a�  �@��ܜ  �Ƀ=��t����$�  �����z�����������������̃��$�m�  �   ��ÍT$��  R��<$�D$tQf�<$t�Ю  �   �u���=�� �C�  �   ����@�  �  �u,��� u%�|$ u��襮  �"��� u�|$ u�%   �t����-`��   �=�� ��  �   �����  ZË�U�����3ŉE�SV3�W��9��u8SS3�GWh��h   S�pp��t�=����Hp��xu
���   9]~"�M�EI8t@;�u�����E+�H;E}@�E�������  ;���  ����  �]�9] u��@�E �5lp3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�/  ��;�t� ��  �P�R���Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5ppSSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w��.  ��;�tj���  ���P����Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�pp��t"SS9]uSS��u�u�u�VS�u �hp�E�V����Y�u�������E�Y�Y  �]�]�9]u��@�E9] u��@�E �u�`�  Y�E���u3��!  ;E ��   SS�MQ�uP�u �~�  ���E�;�tԋ5dpSS�uP�u�u�։E�;�u3��   ~=���w8��=   w��-  ��;�t����  ���P�z���Y;�t	� ��  �����3�;�t��u�SW�~������u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��ͬ  ���u������#u�W�����Y��u�u�u�u�u�u�dp��9]�t	�u��l���Y�E�;�t9EtP�Y���Y�ƍe�_^[�M�3�������Ë�U����u�M������u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap�����(  �ȋAl;��t����Qpu�  ���   Ë�U����u�M��'����E����   ~�E�Pj�u��  ������   �M�H���}� t�M��ap��Ë�U��=� u�E����A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u� �  ������   �M�H���}� t�M��ap��Ë�U��=� u�E����A��]�j �u����YY]Ë�U����u�M��)����E����   ~�E�Pj�u聬  ������   �M�H���}� t�M��ap��Ë�U��=� u�E����A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Ph�   �u���  ������   �M�H%�   �}� t�M��ap��Ë�U��=� u�E����A%�   ]�j �u�~���YY]Ë�U����u�M��$����E����   ~�E�Pj�u�|�  ������   �M�H���}� t�M��ap��Ë�U��=� u�E����A��]�j �u����YY]Ë�U���L��3ŉE�S3�V�uW�]ԉ]�]��]؉]܉u��]�9^�  �F9u P�F0h  P�E�SP�ג  ������  j�  j��  W�E��  jW�E��  jW�E��  jh  �E��  ��$�E�9]��|  9]��s  ;��k  9]��b  9]��Y  �Eԉ3��M܈@=   |�E�P�v�tp���/  �}��%  �E���E�~-8]�t(�E�:�t�x�����M�� �G;�~�@@8X�uۋE�SS�v   Ph   �u܉E�jS�A�  �� ����  �M��E�S�v��   W���   QW@Ph   �vS������$����  �E�S�v�   WP�E�W@Ph   �vS�U�����$���`  �E�}����   3҃}�f��U؉Mč��   �_�Z��M����   �MȈ~S8]�tN�M�M�:�tB�I���;ʉM�'��H   ��M��E� �  f�AA�M̋M��	9M�~�M�AA�M�8Y�u�h�   ��   QP�]���j��   PW�N����E�j��   QP�<������   ��$;�tKP�p��u@���   -�   P�������   ��   +�P�������   +�P�������   �z������E��    ���   �E����   �Eĉ��   �E����   �Eȉ��   �EЉ��   �u��3���Y���m�u��&����u������u������u�����3ۃ�C�ˍ��   �;�tP�p����   ǆ�   ��ǆ�   ��ǆ�    �ǆ�      3��M�_^3�[�6������|"  �ȋAl;��t����Qpu�r  �@��V"  �ȋAl;��t����Qpu�L  ��Ë�U��VW3��u�������Y��u'9 �vV�p���  ; �v��������uʋ�_^]Ë�U��VW3�j �u�u蕩  ������u'9 �vV�p���  ; �v��������uË�_^]Ë�U��VW3��u�u�i�  ��YY��u,9Et'9 �vV�p���  ; �v��������u���_^]Ë�U��VW3��u�u�u�3�  ������u,9Et'9 �vV�p���  ; �v��������u���_^]��̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U���(  ��3ŉE����Vtj
�n�  Y��  ��tj��  Y�����   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P�v�������������(�����0���j ǅ����  @��������,����<p��(���P�8pj�~  ̋�U��M����U#U��#�ʉ��]�Pd�5    �D$+d$SVW�(���3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(���3�P�e��u��E������E�d�    ËM�d�    Y__^[��]QË�U��SV�u���   3�W;�to=��th���   ;�t^9uZ���   ;�t9uP�������   �0�  YY���   ;�t9uP�������   � �  YY���   �z������   �o���YY���   ;�tD9u@���   -�   P�N������   ��   +�P�;������   +�P�-������   �"��������   �=��t9��   uP�m�  �7�����YY�~P�E   ����t�;�t9uP�����Y9_�t�G;�t9uP����Y���Mu�V����Y_^[]Ë�U��SV�5pW�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{���t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5pW�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{���t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�V���t��t;�tWj6Y���  P����Y_^Å�t7��t3V�0;�t(W�8����Y��tV�����> Yu����tV�3���Y��^�3��jh���<  ��  �����Fpt"�~l t��  �pl��uj �x  Y����<  �j�1  Y�e� �Fl�=���i����E��E������   ��j�0  Y�u�á���H�D��H�H����   ������   ������   ������   ������   ����3�Ë�U��SW�}3�;�~,V�u���6�u�u�
�  ����tSSSSS�s�����Ou�^_[]Ë�U��SVW�}h�   3�SW�����u�����u3���   <.u4�F8t-jP���   jP�m�  ����tSSSSS���������   ��h�V�]���  ;��   �} �<0�u��@��   ��.��   PVj@�u�;�}u��@sw��_trP�EVj@��@��}u`��s[��t��,uRP�EVj��P�ֳ  ����t3�PPPPP�v�������,�'����������E�wh�V�X�  ��YY�X������_^[]Ë�U��SV�uV�u�u�������3ۅ�tSSSSS�������F@8tPh�j�u�u�Q��������   8^[tPh zj�u�u�/�����]Ë�U���S3�ChU  �]������Y�E���U  W�x� ��]��^�CH�0�E�h��5L�jhQ  W������E���E��E�L�h�hQ  W��  ����t3�PPPPP�K������sX�E��0�  YY��t�e� �E��E��E����0�CH�0�E�E�h��0jhQ  W�Z������}�|�|��}� uI�FP�p��tP�Ӆ�u	�vP�~���Y�FT��tP�Ӆ�u	�vT�g���Y�E�fT �fL �FP�~H���N�u��I����FP�=p3�Y;�tP�ׅ�u	�vP�*���Y�FT;�tP�ׅ�u	�vT����Y�Fh�^T�^L�^P�^H_[�Ë�U���   ��3ŉE��ESV�uW�}��d����E��\�����`����  �   �H(��T����H,�X �   ��X�����h�������  ��d��� ��  �} ��  �>CuW�~ uQhl��u��d����|�����3���tVVVVV������;�t3�f�f�Gf�G��`���;�t�0��d����G  V�������   Y��P���;�s,V��h����  YY����   V��X����  YY����   ��L��� ��l���VP����YY����   ��l���PSP�ɶ  ������   �C��T������l���PW��h����������> t
��P���;�r��L�����r@PVW��X�����  ����t3�VVVVV�������3�9�\���tjS��\���������9�`���tj��T�����`�����������h����u��d�����������tVVVVV�@�������h����3��M�_^3�[�R����Ë�U����  ��3ŉE�SW���  �u����h���P��P���Ph�   ��x���PS���  ��������u3��  �E���0�sH��x���P��
  YY���x  ��x���P������P��t��������YY��p�����t��CH�M��\����D���k���l���� ��X����1jP��d�����<���P�_����F��x���Q��t�����L�����p��������QP���������t3�PPPPP��������p�����l������CH��P����j��P���P��d�����������}��   ��h�����t��� �F�G$�O ��d����ǋV;t6���t������d�����D����P�H��D�������t�����d���|��"��t�����t�ǋ��P�W���d����H��t���uhj�v��x����vPjh��jj ��  �� ��t93���  f!�Ex���@��r�h�   �5����x���P裵  �����@�G��g �F��G���   �}u	��h����F�Ek�V��H�Y��t1��\�����p����CH�K�����X���Y��l������L����F������\�����t-�E�����<0�7�p��u�7�����sT������cL YY�M��p��������    �1�CH�M�_3�[�P����Ë�U���   ��3ŉE��ESV3ۋ�W��h���;�t;�tP�����Y��  ���D0H��  ǅp���   ��t���;���  �9L�0  �yC�&  �y_�  ��h�W���  ��YY����   +ǉ�p�����   �;;��   ǅl���   �L����p���PW�6�f�������u�6�����Y9�p���t��l�������|�~�Ch�S�+�  ��3�YY;�u	�;;��   ��l���QWS��x���h�   P�B�  ����tVVVVV���������l�����h�����x���Ƅ=x��� ����Y��t��t�����? t
G�? � ���3�9�t�����   ��h����u3��vSSSh�   ��x���PQ�"�����;�tZ�~H��t3�7��x���P�  YY��tS��x����%���Y��u!�p������t���C����~�3�9�p���u9�t���t�D����M�_^3�[�5�����jhؽ�R1  3ۉ]��}v�  �    SSSSS������3��,  �E  ���u��N����Np�]�jh�   �8���YY���}�;���   j��%  Y�E�   �Nl�������]��   �u�M���P���Y�E�;���   9]th���u�  YY��t
��   j�%  Y�E�   �^l���y���W����Y�Fpu2���u)�;����W���j�����Ph,�������������e� �   �-�}܋u�3�j�V$  YËu�j�J$  Y��W�K���W�m���YY�E������   �E��<0  Ëu�fp��jh���/  3��u�3��];���;�u�  �    VVVVV������3��{3��};���;�t�3�f97��;�t��h�  �E;�u�M  �    �ɉu�f93u �8  �    j��E�Ph��i�  ���P�uWS�m�  ���E��E������	   �E��x/  ��u� @  YË�U���SV�u3ۉ]�;�t9]u3��{  v3�f�W�};�u�  SSSSS�    �������<  �u�M�膸���E�;���   9XuH9]v�M��9f�f�8tAFF�M�;Mr�8]�t�E�`p��E���   8]�t�E�`p�����   �uVj�W�=lpj	�p��;���   �Hp��zt�  � *   3�f��   �E�u�E�;�t'��M�:�t�M���QP�w�  YY��tF8t!F9]�u��u+u�u�E�V�uj�p��;�uT�  �M� *   3�f��-9Xu	W�����Y�1SSj�Wj	�p�lp;�u�u  � *   8]�t�E�`p�����H8]�t�M�ap�_^[�Ë�U���SV�u3ۉ]�;�u9]t*�9]w�%  j^SSSSS�0�"���������   3�f�W�};�t��u�M������E;Ev�E=���v	��  j�P�M�QP�uV����������u;�t3�f��  � 8]�tk�M�ap��b@;�tH;Ev<�}�t,3�f��  j"^SSSSS�0������8]�t�E�`p����&�E�E�P   3�f�LF�;�t�8]�t�E�`p��E�_^[�Ë�U��j �u�u�u�u�u�������]�������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[�jh0��v+  j�v   Y�e� �u�N��t/�����E��t9u,�H�JP����Y�v����Y�f �E������
   �e+  Ë���j�A  Y��̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�2���3��ȋ��~�~�~����~���������F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  ��3ŉE�SW������P�v�tp�   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R�o�����C�C��u�j �v�������vPW������Pjj ��  3�S�v������WPW������PW�vS�C�����DS�v������WPW������Ph   �vS������$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[�9�����jhP��V(  �s  ������Gpt�l t�wh��uj �(d  Y���n(  �j�(  Y�e� �wh�u�;5��t6��tV�p��u����tV�D���Y����Gh�5���u�V�p�E������   뎋u�j��  YË�U���S3�S�M��a��������u��   �|p8]�tE�M��ap��<���u��   �xp�ۃ��u�E��@��   ��8]�t�E��`p���[�Ë�U��� ��3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�����   �E��0=�   r����  �p  ����  �d  ��P��p���R  �E�PW�tp���3  h  �CVP菳��3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�H����M��k�0�u��� ��u��*�F��t(�>����E�����D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C����Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95��X�������M�_^3�[�4�����jhp��Q%  �M���j  ���}�������_h�u�u����E;C�W  h   �
���Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�p��u�Fh=��tP� ���Y�^hS�=p���Fp��   �����   j�  Y�e� �C� ��C�$��C�(�3��E��}f�LCf�E�@��3��E�=  }�L����@��3��E�=   }��  ����@���5���p��u���=��tP�g���Y���S���E������   �0j�"  Y��%���u ����tS�1���Y�  �    ��e� �E��	$  Ã=�� uj��V���Y���   3�Ë�U��V�5���5�p�օ�t!������tP�5�����Ѕ�t���  �'�,�V��p��uV�_  Y��th�P��p��t�u�ЉE�E^]�j ����YË�U��V�5���5�p�օ�t!������tP�5�����Ѕ�t���  �'�,�V��p��uV�^  Y��thH�P��p��t�u�ЉE�E^]���p� ��V�5����p����u�5P��e���Y��V�5����p��^á�����tP�5X��;���Y�Ѓ���������tP��p�����  jh���2"  �,�V��p��uV��]  Y�E�u�F\�3�G�~��t$h�P��p�Ӊ��  hH��u��Ӊ��  �~pƆ�   CƆK  C�Fh��j��  Y�e� �vh�p�E������>   j�  Y�}��E�Fl��u����Fl�vl�+���Y�E������   �!  �3�G�uj�  Y�j�  YË�VW�Hp�5���������Ћ���uNh  j�^�����YY��t:V�5���5T������Y�Ѕ�tj V�����YY�Xp�N���	V�@���Y3�W��p_��^Ë�V��������uj��\  Y��^�jh���   �u����   �F$��tP����Y�F,��tP����Y�F4��tP�׶��Y�F<��tP�ɶ��Y�F@��tP軶��Y�FD��tP譶��Y�FH��tP蟶��Y�F\=�tP莶��Yj�:  Y�e� �~h��tW�p��u����tW�a���Y�E������W   j�  Y�E�   �~l��t#W����Y;=��t����t�? uW�)���Y�E������   V�	���Y��  � �uj��  YËuj��  YË�U��=���tK�} u'V�5���5�p�օ�t�5���5�����ЉE^j �5���5T�����Y���u�x���������t	j P��p]Ë�VW�,�V��p��uV��Z  Y�����^  �5�phx�W��hl�W�L���h`�W�P���hX�W�T��փ=L� �5�p�X�t�=P� t�=T� t��u$��p�P���p�L��<�5T��X���p��������   �5P�P�օ���   ��\  �5L������5P��L������5T��P������5X��T��u������X��  ��teh�>�5L������Y�У�����tHh  j������YY��t4V�5���5T�����Y�Ѕ�tj V�y���YY�Xp�N��3�@��$���3�_^Ë�U��3�9Ev�M�9 t@A;Er�]Ë�U��E3�;���tA��-r�H��wjX]Ë���]�D���jY;��#���]��������u�H�Ã���������u�L�Ã�Ë�U��V������MQ�����Y�������0^]���Q�L$+ȃ����Y銺  Q�L$+ȃ����Y�t�  ��U���(  �h��d��`��\��5X��=T�f���f�t�f�P�f�L�f�%H�f�-D���x��E �l��E�p��E�|����������  �p��l��`�	 ��d�   �����������������@p���j��  Yj �<ph���8p�=�� uj�  Yh	 ��4pP�0p��U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh���  �e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E���  Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[�������3�Ë�U���V�u�M�輣���u�P��  ��e�F�P������Yu��P���  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M��I����E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�:�  �M��E��M��H��EP�ɸ  �E�M����Ë�U��j �u�u�u������]Ë�V����tV����@PV�V肦����^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M�������3�;�u+�	���j_VVVVV�8�������}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�����j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h��SV������3ۅ�tSSSSS�������N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F���t�90uj�APQ��������}� t�E��`p�3�_^[�Ë�U���,��3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�ܸ  3ۃ�;�u�~���SSSSS�0�~��������o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q���  ��;�t���u�E�SP�u��V�u��������M�_^3�[������Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   蚟��9}}�}�u;�u+����j^WWWWW�0葫�����}� t�E�`p����  9}vЋE��� 9Ew	�V���j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�߲  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� 觷  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �S�  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�k�����u�E�8 u���} �4����$�p���WF�߶  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP躵  0�F�U�����;�u��|��drj jdRP蔵  0��U�F����;�u��|��
rj j
RP�n�  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N�.�����u-�3���j^�03�PPPPP�.������}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V襞�����}� t�E��`p�3�_^[�Ë�U���,��3ŉE��ESVW�}j^V�M�Q�M�Q�p�0肳  3ۃ�;�u�$���SSSSS�0�$��������Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P谱  ��;�t���u�E�SV�u���`������M�_^3�[躝���Ë�U���0��3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�ǲ  3ۃ�;�u�i���SSSSS�8�i��������   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW���  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[������Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3���P��6������Y���(r�_^Ë�Vh   h   3�V���  ����tVVVVV蠣����^Ë�U�������]�����]��E��u��M��m��]����]�����z3�@��3���hċ��p��th��P��p��tj �������U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]Ã%  Ë�U��3�9Ej ��h   P��p�����u]�3�@��
]Ã=�
uWS3�9�
W�=Lp~3V�5�
��h �  j �v���p�6j �5���׃�C;�
|�^�5�
j �5����_[�5����p�%�� Ë�VW3�����<���u�����8h�  �0���{�  YY��tF��$|�3�@_^Ã$��� 3����S�$pV���W�>��t�~tW��W�X����& Y������|ܾ��_���t	�~uP�Ӄ�����|�^[Ë�U��E�4ŀ��,p]�jh ��  3�G�}�3�9��u�V  j��T  h�   ��G  YY�u�4���9t���nj�\���Y��;�u�(����    3��Qj
�Y   Y�]�9u,h�  W�r�  YY��uW膡��Y������    �]���>�W�k���Y�E������	   �E��H  �j
�(���YË�U��EV�4ŀ��> uP�"���Y��uj��F  Y�6�(p^]Ë�U���
��
k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �������   ��
�5�ph @  ��H� �  SQ�֋�
����   ���	P����@��
����    ����@�HC����H�yC u	�`�����x�ueSj �p�֡���pj �5���Lp��
���k���
+ȍL�Q�HQP襕���E����
;��v�m��
��
�E����=�
[_^�á�
V�5�
W3�;�u4��k�P�5�
W�5����p;�u3��x��
�5�
��
k�5�
h�A  j�5���`p�F;�t�jh    h   W��p�F;�u�vW�5���Lp뛃N��>�~��
�F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W��p��u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U�����
�Mk��
������M���SI�� VW}�����M���������3���U���
����S�;#U�#��u
���];�r�;�u��
��S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1��
�	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t��
�C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;��u�M�;�
u�%�� �M���B_^[����h�_d�5    �D$�l$�l$+�SVW��1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s35�W��E� �E�   �{���t�N�38�<����N�F�38�,����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t����  �E���|@G�E��؃��u΀}� t$����t�N�38蹋���N�V�3:詋���E�_^[��]��E�    �ɋM�9csm�u)�=Ћ t hЋ�ӣ  ����t�UjR�Ћ���M賛  �E9Xth�W�Ӌ�趛  �E�M��H����t�N�38�&����N�V�3:�����E��H���I�  �����9S�R���h�W���a�  ������U��V�EP��訏���؋��^]� �؋�@�����U��V���؋�-����EtV�u��Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR����YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =MOC�t=csm�u+�h������    ��  �W������    ~�I����   �3�]�jh ������}�]��   �s��s�u������   � �e� ;ute���~;w|��  �����Oȋ1�u��E�   �y t�sh  S�O�t��  �e� ��u��-���YËe�e� �}�]�u��u���E������   ;ut�V  �s����Ë]�u��s������    ~�e����   �Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�'���3�A��  ���3��jhH�������M��t*�9csm�u"�A��t�@��t�e� P�q�Ӓ���E�����������3�8E��Ëe��G
  ̋�U��M�V�uƃy |�Q�I�42���^]Ë�U�����u
�X
  �
  �e� �? �E� ~SSV�E�@�@��p��~3�E����E�M�q�P�GE�P�_�������u
K�������E��E��E�;|�^[�E���j��h�����������    t��	  �e� �	  �M���q	  ������Mj j ���   輐���j,h�������ً}�u�]�e� �G��E��v�E�P�I���YY�E��������   �E��������   �E��������   �x����M���   �e� 3�@�E�E��u�uS�uW藔�����E�e� �o�E������Ëe��5�����   �u�}�~�   �O��O�^�e� �E�;Fsk�ËP;�~@;H;�F�L�QVj W�������e� �e� �u�E������E    �   �E��������E�맋}�u�E܉G��u�蕓��Y�����Mԉ��   �����MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v����Y��t�uV�%���YY�jh�����3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w觞  YY����   SV薞  YY����   �G��M��QP�����YY���   �}�E�p�tH�_�  YY����   SV�N�  YY����   �w�E�pV�8��������   ���t|��W�9Wu8��  YY��taSV��  YY��tT�w��W�E�p�_���YYPV�������9�ڝ  YY��t)SV�͝  YY��t�w违  Y��t�j X��@�E���  �E������E��3�@Ëe��F  3�������jh������E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS�N�����FP�w����YYP�vS�4����E������Z����3�@Ëe��  ̋�U��} t�uSV�u�V������}  �uuV��u �����7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP�|���]Ë�U��QQV�u�>  ���   W�������    t?�������   �0���9t+�>MOC�t#�u$�u �u�u�u�uV����������   �}� u�  �u�E�P�E�PV�u W�^������E���;E�s[S;7|G;wB�G�O����H��t�y u*�X��@u"�u$�u�u j �u�u�u�u�����u���E��E���;E�r�[_^�Ë�U���,�MS�]�C=�   VW�E� �I��I����M�|;�|�]  �u�csm�9>��  �~� ��  �F;�t=!�t="���   �~ ��   �G������    ��  �5������   �u�'������   jV�E��  YY��u��  9>u&�~u �F;�t=!�t="�u�~ u�  ��������    t|��������   ������u3����   ����Y��uO3�9~�G�Lh����}����uF��;7|��	  j�u�d���YYh���M��7���h$��E�P�D����u�csm�9>��  �~�~  �F;�t=!�t="��e  �}� ��   �E�P�E�P�u��u W�6��������E�;E���   �E�9��   ;G|�G�E�G�E��~l�F�@�X� �E��~#�v�P�u�E����������u�M��9E���M�E��}� ��(�u$�]��u �E��u��u�u�uV�u�K����u���E����]����}�} t
jV�:���YY�}� ��   �%���=!���   �����   V����Y����   ���������������   � ����}$ �M���   Vu�u��u$�ۉ���uj�V�u�u�������v�����]�{ v&�} �)����u$�u �u�S�u�u�uV������� �������    t�T  _^[�Ë�U��V�u���F����؋��^]� ��U��SVW�V�����   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������� 3�@_^[]�jh`��O����l����@x��t�e� ���3�@Ëe��E������ӯ���h�����?����@|��t������jh�������5�������Y��t�e� ���3�@Ëe��E������}����hn�(���Y����������U���SQ�E���E��EU�u�M�m�詗  VW��_^��]�MU���   u�   Q臗  ]Y[�� ���á�
Vj^��u�   �;�}�ƣ�
jP�y���YY�����ujV�5�
�`���YY�����ujX^�3ҹ��������� ����P�|�j�^3ҹ��W������������������t;�t��u�1�� B��@�|�_3�^��Ϗ���=� t��  �5������YË�U��V�u���;�r"��0�w��+�����Q�z����N �  Y�
�� V�(p^]Ë�U��E��}��P�M����E�H �  Y]ËE�� P�(p]Ë�U��E���;�r=0�w�`���+�����P�*���Y]Ã� P�,p]Ë�U��M���E}�`�����Q�����Y]Ã� P�,p]Ë�U��V�uW3�;�u�o���WWWWW�    �k�������   �F����   �@��   �t�� �F��   ���F�  u	V�  Y��F��v�vV�W  YP�ڛ  ���F;���   �����   �F�uOV�-  Y���t.V�!  Y���t"V�  ��V�<����  ��Y��Y��P��@$�<�u�N    �~   u�F�t�   u�F   ��N�A���������	F�~���_^]�jTh������3��}��E�P��p�E�����j@j ^V虪��YY;��  ����5����   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@�����   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M��������� ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=��|���=���e� ��~m�E����tV���tQ��tK�uQ��p��t<�u���������4����E� ���Fh�  �FP�O�  YY����   �F�E�C�E�9}�|�3ۋ���5������t���t�N��r�F���uj�X�
��H������P��p�����tC��t?W��p��t4�>%�   ��u�N@�	��u�Nh�  �FP蹏  YY��t7�F�
�N@�����C���g����5����p3��3�@Ëe��E������������Ë�VW����>��t1��   �� t
�GP�$p���@   ;�r��6�W����& Y������|�_^Ë�U��EV3�;�u����VVVVV�    蟀���������@^]Ë�U��QV�uV�����E�FY��u�e���� 	   �N ����/  �@t�J���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,������� ;�t�������@;�u�u�Z�  Y��uV��   Y�F  W��   �F�>�H��N+�I;��N~WP�u�  ���E��M�� �F����y�M���t���t���������������P��@ tjSSQ軘  #����t%�F�M��3�GW�EP�u�  ���E�9}�t	�N �����E%�   _[^�Ë�U�����h   �4���Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U���  贆  ��3ŉE��EV3���4�����8�����0���9uu3���  ;�u'�����0����VVVVV�    �~��������  SW�}�����4��������ǊX$�����(�����'�����t��u0�M����u&�<���3��0� ���VVVVV�    �~�����C  �@ tjj j �u�Ė  ���u�W�  Y����  ��D���  �+����@l3�9H�������P��4�� �����p���`  3�9� ���t���P  ��p��4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P��  Y��t:��4���+�M3�@;���  j��@���SP蠙  �������  C��D����jS��@���P�|�  �������  3�PPj�M�Qj��@���QP�����C��D����hp�����\  j ��<���PV�E�P��(���� �4��p���)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4��p����  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@���艖  Yf;�@����h  ��8����� ��� t)jXP��@����\�  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4��p���B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4��p���b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �hp��;���   j ��,���P��+�P��5����P��(���� �4��p��t�,���;����Hp��@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0��p��t��,�����@��� ��8�����Hp��@�����8��� ul��@��� t-j^9�@���u����� 	   �����0�?��@�������Y�1��(�����D@t��4����8u3��$������    ������  ������8���+�0���_[�M�3�^�n����jh��������E���u�����  ����� 	   ����   3�;�|;��r!�v����8�\���� 	   WWWWW�Xw�����ɋ���������������L1��t�P�g�  Y�}���D0t�u�u�u�.������E�������� 	   �����8�M���E������	   �E��T�����u豕  Y�jh��������E���u����� 	   ����   3�;�|;��r����� 	   SSSSS�v�����Ћ����<�����������L��t�P蚔  Y�]���Dt1�u��  YP��p��u�Hp�E���]�9]�t�.����M������ 	   �M���E������	   �E��s�����u�Д  YË�U��V�u�F��t�t�v�Zv���f����3�Y��F�F^]Ë�U��   �}  ��3ŉE�SV�uWV�������3�9FY������}�FjPPS�ʎ  ������������������|��s
������  ����������������� ��ÊH$����F  ������u�F�������+�ʋǋ��  ��V��+��V���������Z  �������  3�9P0�  �����9Vu�������������<  R�p,�p(���������  ��������� Ã���;p(�0���;x,�'���j ������Qh   ������Q�0��p������j ������������������蘍  ����������������������������;��������������t7������K;�s+���u�J�;�s�H�9
u������� ��@��uЍ�����+�3����L  �@�t�V��:
u������B;�r������������u�������  ��x������    �$����F��   �V��u!�������   +N��@�����   jj j ������蕌  ��;�����u$;�����u�F�8��8
uG@;�r��F    �Yj �������������������M�  �����������������   ;�w�N��t
����   t�~������� �DtG������u��)����������� ������uѭ����������3������������M�_^3�[�}i����jh ������u�����Y�e� �u����Y�E��U��E������   �E��U�������u�4���YË�U��V�uV��  Y���u����� 	   ����MW�uj �uP��p�����u�Hp�3���tP�����Y�����������������D0� ���_^]�jh �������E���u覾���  苾��� 	   ����   3�;�|;��r!�}����8�c���� 	   WWWWW�_q�����ɋ���������������L1��t�P�n�  Y�}���D0t�u�u�u��������E��� ���� 	   �����8�M���E������	   �E��[�����u踏  YË�U���SW�}3�;�u 踽��SSSSS�    �p��������f  W�����9_Y�E�}�_jSP�������;ÉE�|ӋW��  u+G�.  ��OV��+�u���tA�U��u������������D2�t��;�s���:
u�E�3�B;�r�9]�u�E���   ��x��	����    �   �G��   �W;�u�]��   �]��u�+�����������E����D0�tyjj �u�������;E�u �G�M��	�8
u�E@;�r��G    �@j �u��u����������}����:�   9Ew�O��t��   t�G�E��D0t�E�E)E��E�M��^_[�Ë�U��V�u�FW��ty�}��t
��t��uh���F��uV�I���EYU3�V�fw���FY��y����F��t�t�   u�F   W�u�uV����YP��  #����t3��褻���    ���_^]�jh@�������u�!���Y�e� �u�u�u�u�:������E��E������	   �E��������u�[���YË�U��V�uWV��  Y���tP�����u	���   u��u�@Dtj�܋  j���Ӌ  YY;�tV�ǋ  YP� p��u
�Hp���3�V�#�  ������������Y�D0 ��tW�޺��Y����3�_^]�jh`�������E���u覺���  苺��� 	   ����   3�;�|;��r!�}����8�c���� 	   WWWWW�_m�����ɋ���������������L1��t�P�n�  Y�}���D0t�u�����Y�E������� 	   �M���E������	   �E��j�����u�ǋ  YË�U��9EuF�jP;Mu+�1���YY���u3�]ËE�    �6�u�7螃�����Q蟔������tՉ�&3�@]Ë�U���EP耎�����EYu��߃�]��Jx	�
�A�
�R�����YË�U��}�t]�Ss��]Ë�U��S�U�������؃��t��P�+���Y��u��[]Ë�U����  ��3ŉE��M�EV3�W�}�������|�����d�����T���ǅ$���^  ��0����������x���;�u 趸��VVVVV�    �k��������5  ;�t��@@SuzP�����Y�P����t���t�ȃ��������������A$u&���t���t�ȃ������������@$�t �1���VVVVV�    �-k��������  �u�������^���ƅc��� ��t�����<������k  ��d�����P����Y��t0��t���VV��t�������YP�k���YYG�P轍��Y��u��  �<%�1  8G�  3���@���ƅ/��� ��X�����L�����l���ƅa��� ƅ`��� ƅj��� ƅS��� ƅb��� ƅs��� ƅk�����(���G���P�6���Y��t��l�����L���k�
�DЉ�l�����   ��N��   ��   ��*tp��F��   ��It��Lut��k����   �O��6u�G�84u��(�������4�����8����m��3u�G�82u���\��dtW��itR��otM��xtH��Xu�A��j����9��ht(��lt��wt��S����"�G�8lt���k�����s������k�����s�����S��� �������j��� ��H���u������0�������������3�2ۉ�D���8�s���u�<Stƅs����<Cuƅs������ ��\�����ntJ��ct��{t��d�����t����}���Y���d�����t����@�����x��������  ��D�����H�����L�����t��l��� ��  ��\�����o�r  �  ��c�
  jdZ;���  �z  ��g~E��it!��n�g  ��j��� ��t����f
  �
  ��\�����x���-�4  ƅ`����1  3ۃ�x���-u��T���� -C�	��x���+u��l�����d�����t����^�����x�����L��� u��l������x����k��l�����l�����tf��x�����T�����X������0���P��|���PCS��T�����$�������������
  ��d�����t����������x�����P�=���Y��u���������   � � ��a���:�x�����   ��l�����l�������   ��d�����t���������T�����x�����a������0���P��|���PCS��T�����$��������������	  ��x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$����{���������	  ��d�����t����������x�����P�6���Y��u���X��� �_  ��x���et��x���E�I  ��l�����l������5  ��T����e��0���P��|���PCS��T�����$��������������  ��d�����t����D�����x�����-u,��T����-��0���P��|���PCS����������  �	��x���+u/��l�����l�����u!�l������d�����t����������x�����x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$������������  ��d�����t����j�����x�����P�ʆ��Y��u���d�����t�����x����U�����X��� YY��  ��j��� ��  ��T�����<��������QP��D���� ��k���HP�5l��j���Y�Ѓ��  ��u��l���ǅL���   ��s��� ~ƅb�����d�����t���W��x�����@�������YY��L��� t��l�����l������3  ��t������x�����x�������  ��\���ctN��\���su��	|	����  �� u2��\���{��  ��a���3ҋȃ�B������L�3˅���  ��j��� ��  ��b��� �~  �� �����P�#k  Y��t��t������������!��������P�����ǅ���?   ���   �� ���P�����P�~  f�������f�FF�  ��p��  �������HH�{  ���������t3�;�x�����  ��c�����j��� �  �����������  ��s��� ~ƅb���G�?^��u
�wƅa����j �E�j P�Y�����>]u	�]F�E� �f��/����^F<-uB��t>���]t7F:�s�����:�w"*������Ћσ��ǳ�����D�GJu�2���ȊЋ��������D��<]u����  ��H�����D���������x���+u'��l���u��t����d�����t����C�����x���j0^9�x����x  ��d�����t���������x���<xtX<XtT��\���xǅX���   t"��L��� t
��l���u��ǅ\���o   �$  ��d�����t���P�����YY��x����  ��d�����t���������L��� ��x���t��l�����l���}��ǅ\���x   ��   �F��D����������@���������t���WP�j���YY9�@�����  ��j��� �  ��<�����\���c��  ��b��� t��D���3�f���  ��D����  ��  ƅk�����x���-u	ƅ`����	��x���+u'��l���u��t����d�����t���������x�����(��� �J  ���  ��\���xte��\���pt\��x���P����Y����   ��\���ou"��x���8��   ��4�����8��������Rj j
��8�����4����<[�������7��x���P����Y��tr��4�����8�����x������������Y��x�����x�����X�����Й����L��� ��4�����8���t��l���t5��d�����t���������x���������d�����t�����x�������YY��`��� ��@�����   ��4�����8����؃� �ى�4�����8�����   ��@�������   ��\���xt;��\���pt2��x���P血��Y����   ��\���ou��x���8}n���,k�
�'��x���P����Y��tR��x����������Y��x�����X�����L��� ��x����|�t��l���t5��d�����t���������x����X�����d�����t�����x�������YY��`��� t�߃�\���Fu��X��� ��X��� �  ��j��� u8��<�����D�����(��� t��4������8����F���k��� t�>�f�>��H�����c���G��H����`<%u
�G�8%u����t�������������G��x�����H���;�ul��P�e  Y��t!��t�����������G��H���;�uG��t�����x����u�?%uD��H����xnu8������	����*��d�����x�������YY�VS��VP����VS�y�������0���u��T����B]��Y��x����u*��<�����u8�c���u�������� t%������ap������� t
������`p���<���[�M�_3�^�jS���Ë�U���VW�u�M��5P���E�u3�;�t�0;�u,�,���WWWWW�    �(\�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�4*  �M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&苧���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9�uh���P������]Ë�U��W��  W�p�u��p���  ��`�  w��t�_]Ë�U����  �u�6  �5��� ��h�   �Ѓ�]Ë�U��h ���p��th��P��p��t�u��]Ë�U���u�����Y�u��p�j蝸��Y�j躷��YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=@� th@��bh  Y��t
�u�@�Y����h�qhxq����YY��uBhʢ�Kt���\q�$tq�c����=�� Yth���
h  Y��tj jj ���3�]�jh������j蹷��Y�e� 3�C9���   ���E���} ��   �5���Q���Y���}؅�tx�5���<���Y���u܉}�u����u�;�rW����9t�;�rJ�6��������������5����������5��������9}�u9E�t�}�}؉E����u܋}��h�q��q�_���Yh�q��q�O���Y�E������   �} u(��j����Y�u�����3�C�} tj�ε��Y������Ë�U��j j�u�������]�jj j ������Ë�V�9�����V�  V�e  V��U��V��  V�Qx  V��+  V�N��V�c���hǝ苝����$���^Ã=�� u�U���V�5��W3���u����   <=tGV���Y�t���u�jGW�~����YY�=����tˋ5��S�BV��~����C�>=Yt1jS��}��YY���tNVSP�M������t3�PPPPP�;U�������> u��5����V���%�� �' ���   3�Y[_^��5���V���%�� ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�Uw  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�pv  Y��t��M�E�F��M��E���Mv  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9��u�њ��h  ��VS����p��5�;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�{����Y;�t)�U��E�P�WV�}�������E���H����5��3�����_^[�Ë�U�� ���SV�5�pW3�3�;�u.�֋�;�t� �   �#�Hp��xu
jX� ��� �����   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5hpSSS+�S��@PWSS�E��։E�;�t/P�>z��Y�E�;�t!SS�u�P�u�WSS�օ�u�u��S��Y�]��]�W��p���\��t;�u���p��;��r���8t
@8u�@8u�+�@P�E���y����Y;�uV��p�E����u�VW�i����V��p��_^[�Ë�V������W��;�s���t�Ѓ�;�r�_^Ë�V� �� �W��;�s���t�Ѓ�;�r�_^Ë�U��QQV���������F  �V\���W�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ����=�����;�}$k��~\�d9 �=�����B߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]Ë�U������e� �e� SW�N�@��  ��;�t��t	�У��`V�E�P�q�u�3u�� q3��Xp3���p3��E�P��p�E�3E�3�;�u�O�@����u������5��։5�^_[�Ë�U���(3�S�]V�uW�}�E��E��E��E��E��E��E��E�9$�t�5������Y��^#�M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E�L���M��]�Q��]���]���Y����  �K���� "   �  �E�H���M��]�Q��E�   �]���]���Y�j  �E�   �E�H���E�@���]���]���"  �M��E�@��r����E�<��׉M��E�<��Z����E�L�놃�tNIt?It0It ��t����   �E�4���E�,���E�L�����E�L��x����E�   ��������   �E�   �E�$���������������   �$����E�<���E�@���E�H���E����E����E���y����E���m����E� ���E�����E�����M����]���]�M��]�Q�E�   ��Y��u賚��� !   �E��_^[�����������"�����.�7�@��%�� �������3�Ë�U��QQSV���  V�5���uw  �EYY�M�ظ�  #�QQ�$f;�uU�v  YY��~-��~��u#�ESQQ�$j�t  ���rVS�)w  �EYY�d�ES�xt���\$�E�$jj�?�u  �]��EY�]�Y����DzVS��v  �E�YY�"�� u��E�S���\$�E�$jj�~t  ��^[�Ë�U��QQS�]VW3�3��}�;���t	G�}���r���w  j��x  Y���4  j��x  Y��u�=���  ���   �A  h���  S�(�W�B������tVVVVV��J����h  �A�Vj �E� ��p��u&h��h�  V�qB������t3�PPPPP�J����V�t��@Y��<v8V��s����;�j�<�hܒ+�QP�.  ����t3�VVVVV�WJ�����3�hؒSW��-  ����tVVVVV�3J�����E��4Ŭ�SW�-  ����tVVVVV�J����h  h��W�>v  ���2j���p��;�t$���tj �E�P�4����6�Fs��YP�6S��p_^[��j�dw  Y��tj�Ww  Y��u�=��uh�   �)���h�   ����YYË�U��E�<�]Ë�U���5<�蔑��Y��t�u��Y��t3�@]�3�]Ë�U��� S3�9]u �V���SSSSS�    �RJ��������   �MV�u;�t!;�u�'���SSSSS�    �#J��������S�����E�;�w�M�W�u�E��u�E�B   �u�u�P�u��aw  ����;�t�M�x�E����E�PS�<���YY��_^[�Ë�U���uj �u�u�u�5�����]Ë�U���   ��3ŉE��ESV�u3ۃ}W��t�����l�����   Sh�   ��|�����Q�u��x����uP�Ѓ  ����;�uj�Hp��z��   SSS�u�u��t���褃  ����p���;�t_3�FVP�np����YY;�tMS��p�����x���W�u�u��t����f�  ����;�tjV�6p��YY��l����;�u!9�x���tW�;I��Y����M�_^3�[�?���ÍN�QWVP�+  ����tSSSSS�aG����9�x���tW��H��Y3��9]u�Sj�D�W�u�uP�f�  ����t�����P�@j��Y��tɊ�
���,0GG��L��|�뱋�U��E�L�]�jh���<���3��]3�;���;�u�����    WWWWW��G��������S�=�
u8j����Y�}�S�/���Y�E�;�t�s���	�u���u��E������%   9}�uSW�5���q����������3��]�u�j�ԥ��Y������U���0���S�ٽ\�����=� t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=� t�#  ��8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����,  �   [�À�8�����=�� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �8������������(�����s4�H��,ǅr���   �0������������ �����v�@�VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�*�  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����D   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Àzuf��\���������?�f�?f��^���٭^����|��剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����|��剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����t����۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-`���p��� ƅp���
��
�t����������l$�l$�D$���   5   �   t��������� u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t�����������l$��������������l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r ����������|$�l$�ɛ�l$������l$��Ã�,��?�$�������,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  �������� �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u��������Ƀ�u�\$0�|$(���l$�-�������l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8����l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w������|$����<$� �|$$�D$$   �D$(�l$(������<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  �������� �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u��������Ƀ�u�\$0�|$(���l$�-�������l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8����l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w������|$����<$� �|$$�D$$   �D$(�l$(������<$�l$$�Q�����0Z�����0Z�������@���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�p  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��P��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��|������������l������   s������t������������d������   v����떋�U�����3ŉE�j�E�Ph  �u�E� �q��u����
�E�P��D��Y�M�3��b*���Ë�U���4��3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5tp�M�QP�֋lp��t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u��$[����YF;�~[�����wS�D6=   w/������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�~H��Y;�t	� ��  ���E���}�9}�t؍6PW�u��|)����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�hp��t`�]��[�hp9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�[Y��YY�E�;�t+WWVPV�u�W�u��;�u�u��Y2��Y�}���}��t�MЉ�u��%��Y�E��e�_^[�M�3��(���Ë�U���S�u�M��z%���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P��8  YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP��  �� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U��QQ��3ŉE��P�SV3�W��;�u:�E�P3�FVh��V�q��t�5P��4�Hp��xu
jX�P���P�����   ;���   ����   �]�9]u��@�E�5lp3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�c}����;�t� ��  �P�	F��Y;�t	� ��  ���؅�ti�?Pj S�'����WS�u�uj�u�օ�t�uPS�u�q�E�S�#���E�Y�u3�9]u��@�E9]u��@�E�u�����Y���u3��G;EtSS�MQ�uP�u��������;�t܉u�u�u�u�u�u�q��;�tV��/��Y�Ǎe�_^[�M�3��<&���Ë�U����u�M��	#���u$�M��u �u�u�u�u�u�������}� t�M��ap���jh�������M3�;�v.j�X3���;E�@u�{���    WWWWW�.����3���   �M��u;�u3�F3ۉ]���wi�=�
uK������u�E;�
w7j詍��Y�}��u试��Y�E��E������_   �]�;�t�uWS�e%����;�uaVj�5���`p��;�uL9=@�t3V�}���Y���r����E;��P����    �E���3��uj�M���Y�;�u�E;�t�    ���K����jh��������]��u�u�C��Y��  �u��uS�*.��Y�  �=�
��  3��}�����  j趌��Y�}�S�ߌ��Y�E�;���   ;5�
wIVSP���������t�]��5V萔��Y�E�;�t'�C�H;�r��PS�u��D��S菌���E�SP赌����9}�uH;�u3�F�u������uVW�5���`p�E�;�t �C�H;�r��PS�u���C��S�u��h������E������.   �}� u1��uF������uVSj �5����p����u�]j����YË}����   9=@�t,V�����Y��������Vy��9}�ul���HpP�y��Y��_����   �1y��9}�th�    �q��uFVSj �5����p����uV9@�t4V�h���Y��t���v�V�X���Y��x���    3��X������x���|�����u��x�����HpP�tx���Y���ҋ�U��MS3�;�v(j�3�X��;Es�x��SSSSS�    �+����3��A�MVW��9]t�u�V���Y��V�u������YY��t;�s+�Vj �S�i"������_^[]Ë�U��E�T��X��\��`�]Ë�U��E���V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5\���q��Y�j h �����3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�~s�����}؅�u����a  �T��T��`�w\���]���������Z�Ã�t<��t+Ht�Vw���    3�PPPPP�P*����뮾\��\���X��X��
�`��`��E�   P�!q���E�Y3��}���   9E�uj����9E�tP�+���Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.����M܋������9M�}�M�k��W\�D�E����p����E������   ��u�wdS�U�Y��]�}؃}� tj 蹇��Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3�裓��Ë�U����HB�PD�M��U���u����Ãe� SW�E��FPj1Q3�C�E�SP�K������FPj2�u��E�SP�6�����FPj3�u��E�SP�!�����FPj4�u��E�SP������P��FPj5�u��E�SP�������FPj6�u��E�SP�����Vj7�u���E�SP�������F Pj*�u��E�SP������P��F$Pj+�u��E�SP������F(Pj,�u��E�SP������F,Pj-�u��E�SP�v�����F0Pj.�u��E�SP�a�����P��F4Pj/�u��E�SP�I�����FPj0�u��E�SP�4�����F8PjD�u��E�SP������F<PjE�u��E�SP�
�����P��F@PjF�u��E�SP�������FDPjG�u��E�SP�������FHPjH�u��E�SP�������FLPjI�u��E�SP������P��FPPjJ�u��E�SP������FTPjK�u��E�SP������FXPjL�u��E�SP�q�����F\PjM�u��E�SP�\�����P��F`PjN�u��E�SP�D�����FdPjO�u��E�SP�/�����FhPj8�u��E�SP������FlPj9�u��E�SP������P��FpPj:�u��E�SP�������FtPj;�u��E�SP�������FxPj<�u��E�SP�������F|Pj=�u��E�SP������P����   Pj>�u��E�SP��������   Pj?�u��E�SP�{�������   Pj@�u�S�E�P�c�������   PjA�u��E�SP�K�����P����   PjB�u��E�SP�0�������   PjC�u��E�SP��������   Pj(�u��E�SP� �������   Pj)�u��E�SP�������P����   Pj�u��E�SP���������   Pj �u��E�SP��������   Ph  �u��E�SP��������   Ph	  �]�S�E�j P�}�����P���_���   [�Ë�U��V�u����  �v�|%���v�t%���v�l%���v�d%���v�\%���v�T%���6�M%���v �E%���v$�=%���v(�5%���v,�-%���v0�%%���v4�%���v�%���v8�%���v<�%����@�v@��$���vD��$���vH��$���vL��$���vP��$���vT��$���vX��$���v\��$���v`�$���vd�$���vh�$���vl�$���vp�$���vt�$���vx�$���v|�$����@���   �t$�����   �i$�����   �^$�����   �S$�����   �H$�����   �=$�����   �2$�����   �'$�����   �$�����   �$�����   �$����,^]Ë�U��SVW�}�  ���t@h�   j�J����YY��u3�@�E��������tV�+���V�#��YY��ǆ�      �����   �;�t�   P�p�73�_^[]Ë�U��V�u��t5�;��tP�j#��Y�F;��tP�X#��Y�v;5��tV�F#��Y^]Ë�U���S�]V3�W�]�u�9su9su�u��u��E���:  j0j��I����YY�};�u3�@�w  ���   jYj��|I��3�Y�E�;�u�u��"��Y�щ09s��   j�UI��Y�E�;�u3�F�u�"���u��"��YY���  �0�u�{>VjW�E�jP�V����E�FPjW�E�jP�A���	E�FPjW�E��E�jP�)�����<E�tV����Y���뎋E�� ����0|��9��0�@�8 u��7��;u���~�����> u������E�����H����u��H�E�3�A��E���t����   �5p��tP�֋��   ��tP�օ�u���   �!�����   �!��YY�E����   �E����   �E���   3�_^[�Ë�U��V�u��t~�F;��tP�Z!��Y�F;��tP�H!��Y�F;��tP�6!��Y�F;��tP�$!��Y�F;��tP�!��Y�F ;��tP� !��Y�v$;5��tV�� ��Y^]Ë�U���SV�uW3��}��u��}�9~u9~u�}��}�����6  j0j�G����YY;�u3�@�u  j�1G��Y�E�;�u	S� ��Y���89~��  j�G��Y�E�;�uS�f ���u��^ ��Y�҉8�v8�CPjV�E�jP�������CPjV�E�jP������CPjV�E�jP�������CPjV�E�jP�������P��CPjV�E�jP�������C PjPV�E�jP������C$PjQV�E�jP������C(PjV�E�j P������P��C)PjVj �E�P�t�����C*PjTV�E�j P�`�����C+PjUV�E�j P�L�����C,PjVV�E�j P�8�����P��C-PjWV�E�j P�!�����C.PjRV�E�j P������C/PjSV�E�j P�������<�t$S����S����u�����u��������Q����C����0|��9��0�@�8 u��#��;u���~�����> u���jY������E�u�   ��	���I�K� �@�M��C3�@3��9}�t�M�����   ;�tP�p���   ;�t#P�p��u���   �P�����   �E��YY�E����   �E����   ���   3�_^[�Ë�U��ES3�VW;�t�};�w�yj��j^�0SSSSS�v�������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u��2j��j"Y����3�_^[]��������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^�Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w�i��j^�0SSSSS���������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x�����#i��j"Y���낋�U��3�S3�@9]|FVW��t>�EÙ+��E���<��7�E�0��X  YY��u
�M���9�}N�u��^;]~�_^3Ʌ���[��]Ë�U�����3ŉE�V���tS�> tNh��V�Z��YY��t=h��V�Z��YY��uj�E�Pj�w�q��t/�u�V��,��Y�M�3�^�^����j�E�Ph  �w�q��u3��׍E�h��P�MZ��YY��u��xp뻋�U��3�f�Mf;���t@@��r�3�@]�3�]Ë�V3��#��,aB<w������,A<w��������tЊ
��u׋�^�3��
B��A|��Z~��a��w@��Ë�U���|��3ŉE�VW�}��c�����ׁƜ   ������jx�E�P�F���%���  PW�q��u!F@�2�E�P�v�UW  YY��uW����Y��t
�N�~�~�F���Ѓ��M�_3�^����� ��U���|��3ŉE�Vjx�E�P�E%�  j   P���q��u3��.�U������9Et�} t�6W�������V���B��Y;�_t�3�@�M�3�^����Ë�U���|��3ŉE�SVW�}��b�����ׁƜ   �y����q��jx�E�P�F���%���  PW�Ӆ�u�f 3�@�b  �E�P�v�@V  YY����   jx�E�P�F���%���  PW�Ӆ�t��E�P�6�V  YY��u�N  �~�R�FuO�F��t,P�E�P�6�%W  ����u�6�N�~�A��Y;Fu!�~��V��uW����Y��t	���V�~�N�   #�;���   jx�E�P�F���%���  PW�Ӆ������E�P�6�eU  Y3�Y��u/�N   �F9^t
   �F�G9^t;�6�}@��Y;Fu.j�9^u49^t/�E�P�6�U  YY��uSW�������YY��t�N   9^u�~�F���Ѓ��M�_^3�[������ ��U���|��3ŉE�VW�}�a�����ׁƜ   ������jx�E�P�F���%���  PW�q��u!F@�[�E�P�6�xT  YY��u	9Fu0j��~ u0�~ t*�E�P�6�RT  YY��uPW���$���YY��t
�N�~�~�F���Ѓ��M�_3�^����� �6�V?���v�����@�F�C?��������f @�~ YY�FtjX���	���jh���F�q�F�   t�   t�u�f ��6��>�������@Y�FtjX������jhb��F�q�Fu�f Ë�U��SVW�_���]���Ɯ   ��u�N  �   �C@�~����t�8 tWjhЛ���������f ��tS�8 tN���t�8 t�������S����~ ��   Vj@hș��������tb�?��t�? t�����P�����I�?��t0�? t+W�>������Y�j@h���F�q�Fu�f ��F  �q�F�F�~ ��   �˃����#ˋ��������}����   ����  ��   ����  ��   ��P��p����   j�v� q����   �E��tf�Nf�f�Nf�Hf�x�]��tm�=q�  f9u%h��j@S�r������t"3�PPPPP������j@Sh  �v�ׅ�t,j@�C@Ph  �v�ׅ�tj
j��S�u�T  ��3�@�3�_^[]Ë�U��VW�}�ǃ� ��  H��  H��  H�I  H��  �M�ESj Z�r  �0;1t|�0�+�t3ۅ��Í\�����i  �p�Y+�t3ۅ��Í\�����H  �p�Y+�t3ۅ��Í\�����'  �p�Y+�t3ۅ��Í\����3����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3����r  �p;qt~�p�Y+�t3ۅ��Í\�����I  �p	�Y	+�t3ۅ��Í\�����(  �p
�Y
+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����w  �p�Y+�t3ۅ��Í\����3����R  �p;qt~�Y�p+�t3ۅ��Í\�����)  �p�Y+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����x  �p�Y+�t3ۅ��Í\�����W  �p�Y+�t3ۅ��Í\����3����2  �p;qt~�p�Y+�t3ۅ��Í\�����	  �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\����3�����   �p;qtr�p�Y+�t3ۅ��Í\����u}�p�Y+�t3ۅ��Í\����u`�p�Y+�t3ۅ��Í\����uC�p�Y+�t3ۅ��Í\����3���u"��+�;�������σ���  �$�������  �P�;Q�tq���Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����3����v����P�;Q�t}���Q�+�t3҅��T�����N����p��Q�+�t3҅��T�����-����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����}����p��Q�+�t3҅��T����3����X����P�;Q�t}���Q�+�t3҅��T�����0����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T�����^����p��Q�+�t3҅��T����3����9����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�to���Q�+�t3҅��T���u6�p��Q�+�t3҅��T���u�p��Q�+�t3҅��T���t����@��I�+�t3Ʌ����L	����3���u3�[�S  �P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����n����p��Q�+�t3҅��T�����M����p��Q�+�t3҅��T�����,����p��Q�+�t3҅��T����3��������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����x����P�;Q�t}���Q�+�t3҅��T�����P����p��Q�+�t3҅��T�����/����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3����Z����P�;Q�t~�Q��p�+�t3҅��T�����1����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����`����p��Q�+�t3҅��T����3����;����I��@�+�� ���3Ʌ����L	���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����b����p��Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����l����P�;Q�t}���Q�+�t3҅��T�����D����p��Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����s����p��Q�+�t3҅��T����3����N����P�;Q�t~�Q��p�+�t3҅��T�����%����Q��p�+�t3҅��T���������Q��p�+�t3҅��T����������Q��p�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T����3����/���f�P�f;Q�������Q��p�+������3҅��T����  �����P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����i����P�;Q�t}���Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����p����p��Q�+�t3҅��T����3����K����P�;Q�t}���Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T�����r����p��Q�+�t3҅��T�����Q����p��Q�+�t3҅��T����3����,����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T�����3����p��Q�+�t3҅��T����3��������p��Q�+������3҅��T���������������M�u��+�t3҅��T�����   �A�V+�t3҅��T�����   �A�V+�t3҅��T�����   �A�N+���   3Ʌ����L	����   �M�u��+�t3҅��T���uh�A�V+�t3҅��T���uK�A�N랋M�u��+�t3҅��T���u �A�N�p����E�M� �	�_���3�_^]�X�J�V�w���������L�+�7�Y���������-���:���~�������������`�l������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U������SV�uW3��E��}�}��}��FFf�> t����at8��rt+��wt�cJ��WWWWW�    �_�����3��S  �  �3ۃM��	�	  �M�3�AFF�f;���  � @  ;��   ����S��   ��   �� ��   ��tVHtG��t1��
t!���u���9}���   �E�   ����   �ˀ   �   ��@��   ��@�   �E�   �   ����   �E����������   �E��}9}�ur�E�   �� �l��TtX��tCHt/��t��������� �  uC��E9}�u:�e������E�   �09}�u%	U��E�   ��� �  u�� �  ��   ��t3���FF�f;������9}���   �FFf�> t�jVh���.E  �����`���j ��X�FFf9t�f�>=�G���FFf9t�jhĜV�PD  ����u��
��   �DjhМV�1D  ����u����   �%jh�V�D  �������������   �FFf�> t�f9>�����h�  �u�ES�uP��B  ����������E����M��H�M�x�8�x�x�H_^[��jh �� e��3�3��}�j�Z��Y�]�3��u�;5�
��   �����9t[� �@��uH� �  uA�F���w�FP�Y��Y����   ����4�V�]u��YY������@�tPV�u��YYF둋��}��h��j8�y!��Y��������9tIh�  � �� P�  YY�����u�4����Y�������� P�(p����<�}�_;�t�g �  �_�_��_�O��E������   ���Fd��Ë}�j�#X��Y�SVW�T$�D$�L$URPQQh��d�5    ��3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�
  �   �C�
  �d�    ��_^[ËL$�A   �   t3�D$�H3�����U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j��	  3�3�3�3�3���U��SVWj j h��Q�i  _^[]�U�l$RQ�t$������]� ��U����u�M��E����E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]�������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �������U��W�}3�������ك��E���8t3�����_�Ë�U���SV�u�M������]�   ;�sT�M胹�   ~�E�PjS������M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P����YY��t�Ej�E��]��E� Y��D��� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�����$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=� u�E�H���w�� ]�j �u�����YY]Ë�U���(��3ŉE�SV�uW�u�}�M��C����E�P3�SSSSW�E�P�E�P��J  �E�E�VP�H@  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[������Ë�U���(��3ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P�5J  �E�E�VP��D  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�9����Ë�U��MSV�u3�W�y;�u�B��j^�0SSSSS���������   9]v݋U;ӈ~���3�@9Ew��A��j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W����@PWV������3�_^[]Ë�U��Q�M�ASVW������  #�% �  �߉E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��E��<  �U����������U��E�����P������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0��3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��O  �uЉC�E։�EԉC�E�P�uV�������$��t3�PPPPP�������M�_�s^��3�[�2����������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�A���YË�U��E�M%����#�V������t1W�}3�;�tVV��W  YY���>��j_VVVVV�8���������_��uP�u��t	�W  ���W  YY3�^]Ë�U��E���]�jh@���[���e� �u�u�$q�E��/�E� � �E�3�=  �����Ëe�}�  �uj��p�e� �E������E��[���������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h`�h�_d�    P��SVW��1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U��3�@�} u3�]��U��SVWUj j hx�u�`  ]_^[��]ËL$�A   �   t2�D$�H�3�����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�d�5    ��3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�u�Q�R9Qu�   �SQ����SQ����L$�K�C�kUQPXY]Y[� ���jh���X��3ۉ]�j�M��Y�]�j_�}�;=�
}W��������9tD� �@�tP����Y���t�E��|(������ P�$p����4����Y����G��E������	   �E��yX���j�YL��YË�U����UV�uj�X�E�U�;�u��:���  ��:��� 	   ����  S3�;�|;5��r'�:����:��SSSSS� 	   ����������Q  ����W�<��������ƊH��u�q:����W:��� 	   �j�����wP�]�;��  ����  9]t7�@$����E���HjYtHu���Шt����U�E�E��   ���Шu!�:�����9���    SSSSS��������4����M;�r�E�u����Y�E�;�u�9���    �9���    ����h  jSS�u�^  ��D(�E���T,���AHtt�I��
tl9]tg��@�M�E�   �D
8]�tN��L%��
tC9]t>��@�M�}��E�   �D%
u$��L&��
t9]t��@�M�E�   �D&
S�M�Q�uP��4��p���{  �M�;��p  ;M�g  �M��D� ���  �}��  ;�t�M�9
u��� ��]�E�É]�E�;���   �M�<��   <t�CA�M�   �E�H;�s�A�8
u
AA�M�
�u�E�m�Ej �E�Pj�E�P��4��p��u
�Hp��uE�}� t?��DHt�}�
t����M��L�%;]�u�}�
t�jj�j��u�  ���}�
t�C�E�9E�G������D� @u����C��+E�}��E���   ����   K���xC�   3�@�����;]�rK�@�� � t����� ���u�^7��� *   �zA;�u��@���AHt$C���Q|	���T%C��u	���T&C+���ؙjRP�u��  ���E�+]���P�uS�u�j h��  �lp�E���u4�HpP�7��Y�M���E�;EtP�X���Y�E�����  �E��  �E��3�;�����E��L0��;�t�M�f�9
u��� ��]�E�É]�E�;���   �E�f����   f��tf�CC@@�E�   �M����;�s�Hf�9
u���Ej
�   �M�   �Ej �E�Pj�E�P��4��p��u
�Hp��u[�}� tU��DHt(f�}�
t�jXf���M��L��M��L%��D&
�*;]�uf�}�
t�jj�j��u�|  ��f�}�
tjXf�CC�E�9E�������t�@u��f� f�CC+]�]������Hpj^;�u�W5��� 	   �_5���0�i�����m�Y����]��\���3�_[^��jh���\R���E���u�'5���  �5��� 	   ����   3�;�|;��r!��4���0��4��� 	   VVVVV��������ɋ���������������L9��t�����;M�Au�4���0�4���    �P��  Y�u���D8t�u�u�u�~������E���`4��� 	   �h4���0�M���E������	   �E��Q����u�  YË�U��QQ�EV�u�E��EWV�E���  ���Y;�u�4��� 	   �ǋ��J�u�M�Q�u�P��p�E�;�u�Hp��t	P��3��Y�ϋ������������D0� ��E��U�_^��jh����P������u܉u��E���u�3���  �3��� 	   �Ƌ���   3�;�|;��r!�r3���8�X3��� 	   WWWWW�T������ȋ���������������L1��u&�13���8�3��� 	   WWWWW������������[P�=  Y�}���D0t�u�u�u�u�������E܉U����2��� 	   ��2���8�M���M���E������   �E܋U��P����u�z  YË�U��E���u�2��� 	   3�]�V3�;�|;��r�b2��VVVVV� 	   �^�����3���ȃ����������D��@^]Ë�U�����3ŉE�V3�95 �tO�=4��u�N  �4����u���  �pV�M�Qj�MQP�0q��ug�= �u��Hp��xuω5 �VVj�E�Pj�EPV�,qP�hp�4����t�V�U�RP�E�PQ�(q��t�f�E�M�3�^������� �   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��"����E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�lp���E�u�M;��   r 8^t���   8]��e����M��ap��Y����0��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�lp���:���뺋�U��j �u�u�u�������]Ë�U��EVW��|Y;��sQ���������<�������<�u5�=��S�]u�� tHtHuSj��Sj��Sj��4q��3�[���/��� 	   ��/���  ���_^]Ë�U��MS3�;�VW|[;��sS������<����������@t5�8�t0�=��u+�tItIuSj��Sj��Sj��4q���3���F/��� 	   �N/������_^[]Ë�U��E���u�2/���  �/��� 	   ���]�V3�;�|";��s�ȃ�����������@u$��.���0��.��VVVVV� 	   ������������ ^]�jh����K���}����������4����E�   3�9^u6j
��@��Y�]�9^uh�  �FP�����YY��u�]��F�E������0   9]�t�������������D8P�(p�E��K���3ۋ}j
�?��YË�U��E�ȃ����������DP�,p]�jh ��"K���M��3��}�j�V?��Y��u����b  j�@��Y�}��}؃�@�<  �4�������   �u�����   ;���   �Fu\�~ u9j
�?��Y3�C�]��~ uh�  �FP�����YY��u�]���F�e� �(   �}� u�^S�(p�FtS�,p��@낋}؋u�j
�>��YÃ}� u��F��+4�����������u�}��uyG�+���j@j �N��YY�E���ta�������� ���   ;�s�@ ���@
�` ��@�E������}�����σ��������DW�����Y��u�M���E������	   �E���I���j��=��Y�����V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U��E���]Ë�U����u�M������E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u�Dp�M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�}  Y����  �t�Etj�c  Y����v  ����   �E��   j�A  �EY�   #�tT=   t7=   t;�ub��M�������{L�H��M�����{,���2��M�����z�����M�����z� ��� ���������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�x  �M��]�� �����������}�E���Hs�S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}�M&��� "   ]��@&��� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3����;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P��������uV�,���Y�E�^�Ë���h��  �u(�  �u�����E ���Ë�U��=� u(�u�E���\$���\$�E�$�uj�/�����$]��)%��h��  �u� !   �J  �EYY]Ë�S��QQ�����U�k�l$���   ��3ŉE��s �CP�s��������u"�e���CP�CP�s�C �sP�E�P�I������s�p������=� u+��t'�s �C���\$���\$�C�$�sP�r�����$�P�����$��  �s �  �CYY�M�3��]�����]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj���  f;�u�E�� u9Utj��3�]Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������"Q���EQQ�$����������  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�-(��]���t����-(��]�������t
�-4��]����t	�������؛�� t���]����jh(��z?��3�9tV�E@tH9@�t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%@� �e��U�E�������e��U�Z?��Ë�U���SVW�����e� �=�� ����   hܤ�8q�����*  �5�phФW�օ��  P����$��W�����P����$��W�����P�����$��W�����P����Y�����thx�W��P����Y������;�tO9��tGP�"���5�������YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9���;�t0P����Y��t%�ЉE���t���;�tP���Y��t�u��ЉE��5�����Y��t�u�u�u�u����3�_^[�Ë�U��MV3�;�|��~��u����(��������> ��VVVVV�    �:��������^]��A@t�y t$�Ix��������QP�zR��YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u����8*u�ϰ?�d����} �^[]Ë�U���x  ��3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������
�����u5����    3�PPPPP�	����������� t
�������`p������
  �F@u^V�Q��Y�P����t���t�ȃ��������������A$u����t���t�ȃ������������@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw�������3��3�3���� �j��Y������;���	  �$�.��������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P����������Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u�H�������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P�8  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  �D�������P����Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7���������5  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V�����������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5h��B��Y�Ћ���������   t 9�����u������PS�5t����Y��YY������gu;�u������PS�5p�����Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�!�����0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u�D��������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF�2  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t����������������� Y���������������t������������������������� t
�������`p��������M�_^3�[�����Ð)&*$Z$�$%%U%�&��U����u�M��ƺ���u�u�u�u�<q�}� t�M��ap��Ë�U��QQ��3ŉE����S�<qVW3�3�G;�u,VVWV�Ӆ�t�=���/�Hp��xu
jX�����������   ;���   ;�u#9uu�E� �@�EVV�u�u�ӋȉM�;�u3��   ~Ej�3�X���r9�D	=   w�M����;�t����  ���P�����Y;�t	� ��  �����3�;�t��u�W�u�u�Ӆ�t VV9uuVV��u�uj�WV�u�hp��W�o���Y����u�u�u�u�q�e�_^[�M�3�膼���Ë�U����u�M��S����u�E��u�u�u�uP�������}� t�M��ap��Ë�S��QQ�����U�k�l$���   ��3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|����G�������uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�������h��  ��x����b����>YYt�=� uV�Q���Y��u�6����Y�M�_3�^������]��[Ë�U��UV�uW��H�F��w�� �
�y�B��w�� ��t;�t�_+�^]Ë�U���S�u�M�蝷��3�9]u.���SSSSS�    ������8]�t�E��`p������   W�};�u+�i��SSSSS�    �e�����8]�t�E��`p������U�E�9XuW�u�:���YY�4V�E� �M�QP�e����E����M�QP�S�����G;�t;�t�+���^8]�t�M��ap�_[�Ë�U��V3�95�u09uu����VVVVV�    ������������9ut�^]����V�u�u�������^]Ë�U���S3�VW9]��   �u�M��i���9]u.�m��SSSSS�    �i�����8]�t�E��`p������   �};�t˾���9uv(�.��SSSSS�    �*�����8]�t�E��`p����`�E�9Xu�uW�u��,  ��8]�tD�M��ap��;�E� �M�QP�����E����M�QP������G�Mt;�t;�t�+����3�_^[�Ë�U��V3�95�u99uu���VVVVV�    �����������'9ut܁}���w�^]�H,  V�u�u�u������^]Ë�U��QSV��3�;�u�3��j^SSSSS�0�0��������   W9]w���j^SSSSS�0���������   3�9]���A9Mw	����j"�ЋM�����"w��]���9]t�-�N�E�   �؋�3��u��	v��W���0�A�E�3�;�v�U9U�rڋE�;Er�럈I���I�G;�r�3�_^[�� ��U��}
�Eu
��}jj
�j �u�u�M�����]Ë�U���4S3��E�VW���]��]��E�   �]�t	�]��E��
�E�   �]��E�P�-  Y��tSSSSS�վ�����M� �  ��u�� @ u9E�t�M������+ú   ��   �tGHt.Ht&����������j^SSSSS�0覿�����  �U����t��   u��E�   @��}��EjY+�t7+�t*+�t+�t��@u�9}����E���E�   ��E�   ��E�   ��]��E�   #¹   ;��   ;t0;�t,;�t=   ��   =   �@����E�   �/�E�   �&�E�   �=   t=   t`;������E�   �E�E�   ��t�����#M��x�E�   �@t�M�   �M�   �M��   t	}�� t�M�   ��E�   릨t�M�   �c�������u�]������@���    �   �E�=@qS�u��    �u�E�P�u��u��u�׉E���um�M��   �#�;�u+�Et%�e����S�u�E��u�P�u��u��u�׉E���u4�6�������������D0� ��HpP��
��Y�
��� �u  �u���p;�uD�6�������������D0� ��Hp��V�
��Y�u�� p;�u��R
���    룃�u�M�@�	��u�M��u��6�������Ѓ�������Y��Y�M����L��Ѓ����������D$� ��M��e�H�M���   �����  �Etrj���W�6�J�����E�;�u��	���8�   tN�6�_N�������j�E�P�6�]���������uf�}�u�E�RP�6��'  ��;�t�SS�6�FJ����;�t��E���0  � @ � @  �}u�E�#�u	M�	E�E#�;�tD=   t)= @ t"=   t)= @ t"=   t= @ u�E���M�  #�;�u	�E���]��E   ��  �E�@�]���  �E��   �#�=   @��   =   �tw;���  �E�;��y  ��v��v0���f  �E�3�H�&  H�R  �E���  �E�   �  jSS�6�*������t�SSS�6����#���������j�E�P�6�?���������t�����tk����   �}�﻿ uY�E���   �E�;���   ���b������P���jSS�6��������C���SSS�6������#����   �����E�%��  =��  u�6�TL��Y���j^�0���d  =��  uSj�6�XH�������������E��ASS�6�=H������E�﻿ �E�   �E�+�P�D=�P�6�B������������9}�ۋ�������������D$�2M���0��������������D$�M�������
ʈ8]�u!�Et��ȃ����������D� �}��   ���#�;�u|�Etv�u�� pS�u�E�jP�u������W�u�@q���u4�HpP�����ȃ����������D� ��6����Y�����6���������������_^[��jhH��P#��3��u�3��};���;�u����j_�8VVVVV����������Y��3�9u��;�t�9ut�E%������@tu��u�u�u�u�E�P���i������E��E������   �E�;�t���	#���3��}9u�t(9u�t��������������D� ��7�=���YË�U��j�u�u�u�u�u������]Ë�U���SV3�3�W9u��   �];�u"���VVVVV�    �����������   �};�t��u�M��ԫ���E�9pu?�f��Ar	f��Zw�� ���f��Ar	f��Zw�� CCGG�M��tBf��t=f;�t��6�E�P�P�%  ���E�P�P�u%  ��CCGG�M��t
f��tf;�t�����+��}� t�M��ap�_^[�Ë�U��V3�W95�u3�9u��   �};�u�#��VVVVV�    �����������`�U;�t��f��Ar	f��Zw�� ���f��Ar	f��Zw�� GGBB�M��t
f;�tf;�t�����+��V�u�u�u�w�����_^]Ë�U��} u3�]ËU�M�Mt�f��tf;uAABB����
+�]Ë�U����  ��f9Eu�e� �e�   f9Es�E���f�Af#E���E��@�u�M������E��p�p�E�Pj�EP�E�jP�$  ����u!E��}� t�E�`p��E��M#��Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5�N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC����+�;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5�N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3���A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ; �����   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}� ����3�@�   ���e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+���M���Ɂ�   �ً�]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5 �N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC����+ �;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5 �N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��$�A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;��$���   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}���,��3�@�   �,��e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+$���M���Ɂ�   �ً(�]���@u�M�U�Y��
�� u�M�_[�Ë�U���|��3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u����SSSSS�    ������3��O  �U�U��< t<	t<
t<uB��0�B���/  �$��P�Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �#  =�����/  �����`�E�;���  }�ع ��E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9U�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �;����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[覛����cJ�JK@K�K�K�K,LL�L�L:L��U���t��3ŉE�S�]VW�u�}�f��E��U�� �  #��E��A�#�f�}� �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   t�C-��C �u�}�f��u1��u-��u)3�f9M�f�����$ �C�C�C0�C 3�@�  f;���   3�@f��   �;�u��t��   @uh���Sf�}� t��   �u��u;h���;�u0��u,h���CjP������3���tVVVVV�������C�*h���CjP�ř����3���tVVVVV�������C3��s  �ʋ�i�M  �������Ck�M��������3���f�M๠��ۃ�`�E�f�U�u�}�M�����  }� ��ۃ�`�E�����  �E�T�˃������h  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��z����M�����?  ��  f;���  �]��E�3��ɉU��U��U�U��U�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��U���3�3�f9u���H%   � ���E��[���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �_�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[茒���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��q���Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��3�PPjPjh   @h���Dq�4�á4�V�5 p���t���tP�֡0����t���tP��^á���3�9������Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v�\���j^SSSSS�0�Y��������V�u�M��-����E�9X��   f�E��   f;�v6;�t;�vWSV�<������	���� *   ������ 8]�t�M��ap�_^[��;�t2;�w,�����j"^SSSSS�0�ە����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�hp;�t9]�^����M;�t����Hp��z�D���;��g���;��_���WSV�e������O�����U��j �u�u�u�u�|�����]�U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U���SVW3�jSS�u�]��]��e����E�#��U���tYjSS�u�I�����#ʃ����tA�u�}+����   ;���   �   Sj�LqP�`p�E���u�2����    �'���� _^[��h �  �u�  YY�E���|
;�r�����P�u��u��������t6�+��xӅ�wϋu��u��u��   YY�u�j �LqP�Lp3��   ������8u�����    ����u��;�q|;�skS�u�u�u�N���#�����D����u�7���YP�Hq�����H��E�#U���u)�F����    �N������Hp��u�#u��������S�u��u��u����#���������3��������U��S�]V�u��������������0�A$�W�y����   ���� @  tP�� �  tB��   t&��   t��   u=�I��
�L1$��⁀���'�I��
�L1$��₀���a��I��
�L1$�!���_^[u� �  ]����% �   @  ]Ë�U��EV3�;�u�.���VVVVV�    �*�����jX�
����3�^]Ë�U����  �ȃ�f9M��   S�u�M��օ���M�Q3�;�u�E�H�f��w�� ���aV�   ��f9u^s)�E�Pj�u�9��������Et9�M싉�   f����q�M�jQj�MQPR�E�P�*  �� ���Et�E�8]�t�M�ap�[�Ë�U����u�M��3����}�}3���u�u�u�u�q�}� t�M��ap��Ë�U�����3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[�Z����Ë�U����u�M��'����E��~�M��Jf�9 t	AA��u���+�H�u �uP�u�u�u�pp�}� t�M��ap����%Pp�����̋T$�B�J�3���������s�������̋T$�B�J�3��ą������S�������̋T$�B�J�3�褅���t��3�������̋T$�B�J�3�脅���̵��������̋T$�B�J�3��d����$���������̋T$�B�J�3��D������ӏ������̋T$�B��h���3��!����J�3������ȷ馏���������̋T$�B�����3������T�透���̋T$�B�J�3��Ԅ���Ը�c�������̋T$�B�J�3�贄���J�3�誄���,��9�������������̋T$�B�J�3�脄�������������̋T$�B�J�3��d����ܹ��������̋T$�B�J�3��D����4��ӎ������̋T$�B�J�3��$����J�3��������驎���M���w���T$�B�J�3��������醎���M���0���T$�B�J�3��ԃ�����c����M��0���M����ҡ���T$�B�J�3�覃���L��5����M��w���u��n��YËT$�B�J�3��y�����������M�邡���T$�B�J�3��V�����������T$�B�J�3��;�������ʍ��������������h`i蒧��Yù ��xv��h�i�|���Y�h�i�p���Yù���Vv��h�i�Z���Y�h�i�N���YÃ=�� uK�����t�t��Q<P�B�Ѓ����    �����tV������V�m�������    ^ù ��v���D��W/�������u������~��                                   �� 
� � *� <� �� �� �� �� �� �� �  � 4� H� d� �� �� �� �� �� �� �� �� � � "� 8� N� ^� j� t� �� �� �� �� �� �� �� �� �� � � *� 8� H� V� h� x� �� �� �� �� �� �� �� �� � � 6� N� h� �� �� �� �� �� �� �� � � 4� J� Z� �� �� �� �� �� �� �� �� � �     f�         i>iTii2i        ?�;:E�n��        D^�o                    ���N       �   p� p� bad allocation  ���! � P ��@ ��� � �o3D-COAT     c:\program files\maxon\cinema 4d r13 demo\plugins\applink_cinema4dr13\source\applinkdialog.cpp  Start import!   To import a new object? File exists!    export.txt  Folder ..\MyDocuments\3D-CoatV3\Exchange not found! 3D-CoatV3   Exchange    preference.ini  3D-Coat.exe is run! 3D-Coat.exe not found!  open                c:\program files\maxon\cinema 4d r13 demo\plugins\applink_cinema4dr13\source\applinkexporter.cpp    
   c:\program files\maxon\cinema 4d r13 demo\resource\_api\ge_dynamicarray.h   ]   autopo  curv    prim    alpha   vox retopo  ref uv  ptex    mv  ppp [   # end   v       # begin      vertices
        �?vt   texture vertices
  /   f   usemtl   faces
 g   mtllib  mtl map_    illum 2
    Tr 0.000000
    Ns 50.000000
   Ks  Kd  Ka 0.300000 0.300000 0.300000
  newmtl  No selected objects!    Object "    " has no UVW tag.
UV coordinates can't be exported. Material not found on   object. Default Name    Export object   #Cinema4D Version:  %d.%m.%Y  %H:%M:%S  #File created:  #Wavefront OBJ Export for 3D-Coat
  File     write success! [SkipExport]
   [SkipImport]
         �import.txt  output.obj  obj x�� ����p� ���� L� � 0��� D��� @�  � �� p� �� ��  � P� @� ��       Y@��`� � �  � 0� �� @� ` � �� � `�  � p� ܪ�� �0�  � �� �� @� ` � �� @� `�  � p� (�p� �� �� �� p� p� �� �� Selection   Error on inserting phongTag. Object:    Create objects...   Memory allocation error for material.   x��
Ы�(�� � 00@� ` � �� ���2���h��������vector<T> too long  bad cast    ios_base::eofbit set    ios_base::failbit set   ios_base::badbit set    T��7    X       P   f   vt  Gathering of data...     not found!  can not removed!   normalmap   displacement %f displacement    map_Ks %s   map_Ks  map_Kd %s   map_Kd  Ke %lf %lf %lf  Ke  Ks %lf %lf %lf  Ks  Ka %lf %lf %lf  Ka  Kd %lf %lf %lf  Kd  illum %d    illum   d %lf   d   Ns %lf  Ns  newmtl %s   Open file   .       c:\program files\maxon\cinema 4d r13 demo\plugins\applink_cinema4dr13\source\applinkimporter.cpp    vt %lf %lf %lf  vt %lf %lf  v %lf %lf %lf   g %s    mtllib %s   Parse file...   Open file:  textures.txt    ��I�H����`�Їp�����icon_coat.tif   c:\program files\maxon\cinema 4d r13 demo\plugins\applink_cinema4dr13\source\applinkpreferences.cpp     c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_file.cpp         �f@-DT�!	@h���������М������o�������������     @�@|���������М������Ȯ��p���� ����0� �@� �c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_gui.cpp ���������М�����0�    \���������М������p�����������к�� �0���Progress Thread 0%  ~   %       c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_general.h   %s     ����MbP?��iPO(��i    c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_baseobject.cpp      c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_resource.cpp    #   M_EDITOR    t� �res c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_pmain.cpp   c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_basetime.cpp              �? �Ngm��C   ����A  4&�k�  4&�kC�� � � ��    c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_libs\lib_ngon.cpp   c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_basebitmap.cpp  а��    c:\program files\maxon\cinema 4d r13 demo\resource\_api\c4d_gv\ge_mtools.cpp    ���`�`��������*   C   ����@����string too long invalid string position r            
   !   "   2   *            #   3   +       w   a   r b     w b     a b     r +     w +     a +     r + b   w + b   a + b   ����+�����ز���Unknown exception   �?���csm�               �                      �?      �?3      3            �      0C       �       ��                                                                                                                                                                                                                                                                                                        ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������LC_TIME LC_NUMERIC  LC_MONETARY LC_CTYPE    LC_COLLATE  LC_ALL  8�    ^#,���^# ���_��������q� �����	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ _., _   ;   =   =;  EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    `���e+000          �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    jc8�ua��bad exception   CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:                �������             ��      �@      �              �?5�h!���>@�������             ��      �@      �        HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun united-states   united-kingdom  trinidad & tobago   south-korea south-africa    south korea south africa    slovak  puerto-rico pr-china    pr china    nz  new-zealand hong-kong   holland great britain   england czech   china   britain america usa us  uk  swiss   swedish-finland spanish-venezuela   spanish-uruguay spanish-puerto rico spanish-peru    spanish-paraguay    spanish-panama  spanish-nicaragua   spanish-modern  spanish-mexican spanish-honduras    spanish-guatemala   spanish-el salvador spanish-ecuador spanish-dominican republic  spanish-costa rica  spanish-colombia    spanish-chile   spanish-bolivia spanish-argentina   portuguese-brazilian    norwegian-nynorsk   norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg   german-lichtenstein german-austrian french-swiss    french-luxembourg   french-canadian french-belgian  english-usa english-us  english-uk  english-trinidad y tobago   english-south africa    english-nz  english-jamaica english-ire english-caribbean   english-can english-belize  english-aus english-american    dutch-belgian   chinese-traditional chinese-singapore   chinese-simplified  chinese-hongkong    chinese chi chh canadian    belgian australian  american-english    american english    american    ��ENU ��ENU ��ENU ��ENA ��NLB t�ENC p�ZHH l�ZHI d�CHS P�ZHH <�CHS (�ZHI �CHT �NLB �ENU �ENA ԘENL ȘENC ��ENB ��ENI ��ENJ ��ENZ t�ENS X�ENT L�ENG @�ENU 4�ENU $�FRB �FRC  �FRL �FRS ��DEA ̗DEC ��DEL ��DES ��ENI ��ITS |�NOR h�NOR T�NON <�PTB (�ESS �ESB �ESL ��ESO ��ESC ĖESD ��ESF ��ESE ��ESG x�ESH h�ESM X�ESN D�ESI 4�ESA  �ESZ �ESR ��ESU �ESY ؕESV ȕSVF ��DES ��ENG ��ENU ��ENU ��USA ��GBR ��CHN ��CZE ��GBR |�GBR t�NLD h�HKG \�NZL X�NZL L�CHN @�CHN 4�PRI ,�SVK �ZAF �KOR  �ZAF ��KOR ��TTO ��GBR ДGBR ��USA ��USA 6-0   OCP ACP Norwegian-Nynorsk   c c s   U T F - 8   U T F - 1 6 L E     U N I C O D E    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   ->* &   +   -   --  ++  ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        p�h�\�P�D�8�,�$����r`�D�0����������������ءԡh�С̡ȡġ�����tH}������������D}������������������|�x�t�p�l�`�T�L�@�(����Ƞ����h�D�(�������������t�P�H�<�,���Ȟ��x�L�0�������t��r_nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    1#QNAN  1#INF   1#IND   1#SNAN  CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           ���   RSDS�����6�I�@(,��   C:\Program Files\MAXON\CINEMA 4D R13 Demo\plugins\Applink_Cinema4DR13\obj\Applink_Cinema4DR13_Win32_Release.pdb             ��           �(�D�    �       ����    @   � �        ����    @   `�           p�D�                @���           ����ħ    @�       ����    @   ��\�        ����    @   �           �ħ                x��           �$�    x�        ����    @   �           P�\�$�    ��       ����    @   @�           ����$�    ��       ����    @   x�            ��Ĩ           Ԩ���    ��       ����    @   Ĩ��       ����    @   �           (�0�    ��        ����    @   �           �`�           p��������    �       ����    @   `�L�              P   ��           ̩ܩ���    L�       ����    @   ����              @   Ĩ��              @   �            L���            ��X�           h�x���$�    ��       ����    @   X�            ����           ����    ��        ����    @   ��            ���            ����    ��       ����    @   �            0�<�           L�\�\�$�    0�       ����    @   <�    P       P���           �����������    P�       ����    @   ��            ���           �� ���    ��       ����    @   �            ��0�           @�L�ħ    ��       ����    @   0�             �|�           ����ħ     �       ����    @   |�             �Ȭ           ج�L�ħ     �       ����    @   Ȭ            @��           (�8���ħ    @�       ����    @   �    X       ��h�           x����������    ��       ����    @   h�           ��ȭ�    ��       ����    @   ����        ����    @    �           ��                ��,�           <�L�ȭ�    ��       ����    @   ,�             �`�            ,���           ����D�    ,�       ����    @   ��            H�ܮ           ���    H�        ����    @   ܮ            d�$�           4�@�D�    d�       ����    @   $�            |�p�           ����@�D�    |�       ����    @   p�           ��į    ��        ����    @   ��            ����           ��    ��        ����    @   ��            ��<�           L�X�į    ��       ����    @   <�            �� �            <���           ����    <�        ����    @   ��            l��           ����    l�        ����    @   �            ��,�           <�D�    ��        ����    @   ,�            ��t�           ����į    ��       ����    @   t�            ����           бر    ��        ����    @   ��            ���           �$�$�    ��       ����    @   �            $�T�           d�t�L�ħ    $�       ����    @   T�            ����           ����    ��        ����    @   ��            \��            d� �           ��ħ    d�       ����    @    �            ��L�           \�h�ħ    ��       ����    @   L�            � � �_ �� � @f `f �f �f �f �f  g 0g Pg pg �g �g �g  h -h Ph ~h �h �h �h                         ��     �   $�@�    @�    ����       ��     \�    ����       X�            �� ����    ����                  \�"�   l�   |�                            �            ,����    ����                  "�   Դ   �                            Ĵ              ��            �	����    ����                  @�"�   P�   `�                            
����    ����                  ��"�   ��   ��                            �����    ����                  �"�    �   �                    0    X�   h���@�     �    ����    (   `#    ��    ����    (   �"    �    ��   ��@�    d�    ����       ��            �&����    ����                  ض"�   �   ��                    p    @�   P�l�@�    @�    ����    (   �'     �    ����    (   �'            �+            �+����    ����    ����    ����    "�   ��   �                              ��            ��            �/            �.����    ����    ����    ����    "�   4�   x�                              $�            �            2����    ����                  ��"�   ��   ��                             7����    ����                  ��"�   �   �                            9����    ����                  P�"�   `�   p�                            �=����    ����                  ��"�   ��   ȹ                            �?����    ����                   �"�   �    �                            �D            �C����    ����    ����    ����    "�   x�   ��                              h�            X�����%h"�   �                       ����Hh"�   �                       ����kh    sh"�   <�                       �����h    �h"�   p�                       �����h"�   ��                           ��    �   ���@�    $�    ����    (   ^�    ����    ����    ����    	�    ����    ����    ����     �    ����    ����    ����    ,�    ����    ����    ����    ��    ����    ����    ����    �        ������    ����    ����    m�    ����    ����    ����    t     ����    ����    ����    X    ����    ����    ����    �    ����    ����    ����        ����    ����    ������    ����    ����    ����    !    ����    ����    ����    �    ����    ����    ����    �"    ����    ����    ����    j/        (/        9/    ����    ����    ����    .0    ����    ����    ����    E4    ����    ����    ����    �7    ����    ����    ����    d;    ����    ����    ����    �=����     >����    ����    ����    �?����    �?����    ����    �����D�D    ����    ����    ����    ^T    ����    ����    ����    c    �b�b����    ����    �����c�c@           �d����    ����                  d�"�   t�   ��                   ����    ����    ����    �e    <eEe����    ����    �����g�g    ����    ����    ����LhPh    ja    4�   @�@�    ��    ����       m    ����    ����    ����%n)n    ����    ����    ����unyn    ����    ����    ����	tt    ����    ����    ����    R~    ����    ����    ����    3    ����    ����    ����    ��    ����    ����    ����    K�    ����    ����    ����    ӆ    ����    ����    ����    <�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    4�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    `�    ����    ����    ������    ����    ����    ����/    ����    ����    ����    -    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    �        �����    ����    ���� #     ����    ����    ����    �<��         X�  p ��         x� Tq                     �� 
� � *� <� �� �� �� �� �� �� �  � 4� H� d� �� �� �� �� �� �� �� �� � � "� 8� N� ^� j� t� �� �� �� �� �� �� �� �� �� � � *� 8� H� V� h� x� �� �� �� �� �� �� �� �� � � 6� N� h� �� �� �� �� �� �� �� � � 4� J� Z� �� �� �� �� �� �� �� �� � �     f�     C CloseHandle EProcess32Next Module32First CProcess32First  � CreateToolhelp32Snapshot  KERNEL32.dll  ShellExecuteExA SHELL32.dll �InterlockedIncrement  �InterlockedDecrement  !Sleep �InitializeCriticalSection � DeleteCriticalSection � EnterCriticalSection  �LeaveCriticalSection  -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent ZRaiseException  �GetLastError  �HeapFree  �RtlUnwind � DeleteFileA �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �LCMapStringA  zWideCharToMultiByte MultiByteToWideChar �LCMapStringW  [GetCPInfo RGetACP  GetOEMCP  �IsValidCodePage �GetModuleHandleW   GetProcAddress  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �SetLastError  �GetModuleHandleA  �HeapCreate  �HeapDestroy WVirtualFree TVirtualAlloc  �HeapReAlloc �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA �WriteFile �GetConsoleCP  �GetConsoleMode  AFlushFileBuffers  hReadFile  �SetFilePointer  ExitProcess �GetModuleFileNameA  JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW �GetEnvironmentStringsW  TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �HeapSize  �GetLocaleInfoA  =GetStringTypeA  @GetStringTypeW  mGetUserDefaultLCID  � EnumSystemLocalesA  �IsValidLocale �InitializeCriticalSectionAndSpinCount �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW �SetStdHandle  �LoadLibraryA  �GetLocaleInfoW   CreateFileW x CreateFileA �SetEndOfFile  #GetProcessHeap              ���N    b�          X� \� `�  � z�   Applink_Cinema4DR13.cdl c4d_main                                                                                                                              �q<�    .?AVApplinkDialog@@ <�    .?AVGeDialog@@  �q�q<�    .?AVbad_alloc@std@@ <�    .?AVexception@std@@ <�    .?AVfacet@locale@std@@  <�    .?AVcodecvt_base@std@@  <�    .?AUctype_base@std@@    <�    .?AVios_base@std@@  <�    .?AV?$_Iosb@H@std@@ <�    .?AV?$basic_istream@DU?$char_traits@D@std@@@std@@   <�    .?AV?$basic_ios@DU?$char_traits@D@std@@@std@@   <�    .?AV?$ctype@D@std@@ <�    .?AV?$basic_streambuf@DU?$char_traits@D@std@@@std@@     <�    .?AV?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    <�    .?AV?$codecvt@DDH@std@@ <�    .?AV?$basic_istringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    <�    .?AV?$basic_filebuf@DU?$char_traits@D@std@@@std@@   <�    .?AVlogic_error@std@@   <�    .?AVruntime_error@std@@ <�    .?AVlength_error@std@@  <�    .?AVfailure@ios_base@std@@  <�    .?AVbad_cast@std@@  <�    .?AV?$basic_ifstream@DU?$char_traits@D@std@@@std@@  �q�q<�    .?AVCommandData@@   <�    .?AVBaseData@@  <�    .?AVApplinkPreferences@@    �q�q�q�q<�    .?AVGeModalDialog@@ <�    .?AVGeUserArea@@    <�    .?AVSubDialog@@ <�    .?AViCustomGui@@    �q�q�q�q�q�q�q�q�q�q<�    .?AVGeSortAndSearch@@   <�    .?AVNeighbor@@  <�    .?AVDisjointNgonMesh@@  �q�q�q�q�q�q�q�q�q<�    .?AVC4DThread@@ �q�q�q�q�q�q<�    .?AVGeToolNode2D@@  <�    .?AVGeToolDynArray@@    <�    .?AVGeToolDynArraySort@@    <�    .?AVGeToolList2D@@  �q�����q<�    .?AV_Locimp@locale@std@@    �q   �q<�    .?AVout_of_range@std@@  �q����������� ���� �(�0�        �q
   Copyright (c) 1992-2004 by P.J. Plauger, licensed by Dinkumware, Ltd. ALL RIGHTS RESERVED.      �q<�    .?AVtype_info@@ N�@���D            u�  s�          �q            fmod         ����D����}�}���}�����sqrt    ����   ��        �q                                                                                                                                                                                                                                                                                                                                                abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     ���  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����    C                                                                                              ��            ��            ��            ��            ��                              ��        ���� �����   ������������                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                          �q<�    .?AVbad_exception@std@@             ��    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����
                                                          ǝ      x   
   ?     ��   T�	   (�
   ��   d�   4�   �   �   ��   ��   L�   �   �   ̏   h�    0�!   8�"   ��x   ��y   t�z   d��   `��   P�       ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      ���4�:�?�E�J�P�V�\�b�~���������ʳ޳���-�2�R�f�~�������Ѵִ��
�"�6�V�[�u�z�����Ƶڵ������>�R�j�~�������¶����"�B�G�a�f�������  ����������������������t�l�`�\�X�T�P�L�H�D�@�<�8�4�0�(����L���������ԓȓē��������	         ��.   ��h�h�h�h�h�h�h�h�h���   .       �                                                                                                                                                                                                                                   �&         H�   L�   <�   @�   p�   h�!   `�   4�   ,�   �   X�   P�    �   ��    ��   �   �   H�   �   @�   8�   0�   (�    �"   �#   �$   �%   �&    �      �      ���������              �       �D        � 0     ���    �p     ����    PST                                                             PDT                                                             `�������        ����           ���5      @   �  �   ����             ������������   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l           �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                                                       �   0040E0t0�0�0�0�01J142]2�2 323F3~3�3�3�3�3�3�3
4.4E4[4e4m67@7N7f7z7�7	8808A8V8c8x8�8�8�8�8�8�899)9=9P9^9s9�9�90:m::�:�:�:;8;e;�;�;�;<\<�<�<�< =2=D=�=~>�>�>�>�>�>f?p?�?�?�?�?      �   080c0v0�0�0�011%191O1d1�14D4_4s4�4�4�4�4�4l5�5�5�5�5I6^6r6�6�6�6�6�697N7p7�78898�8�89y9�9�9�9
::):p:�:�:�:�:�:�:�:@;�;�;�;<<$<<<g<�<�<�<�<�<==5=M=o=�=�=�=�=�=
>>.>6>I>a>�>�>�>�>�>�>�>�>�>�>�> 0  H  �1�1�1�12"2Z2l2}2�2�2�2�2 333,3>3G3Y3k3s3�3�3�3�3�34(4G4^4s4�4�4�4�4�45!555Q5c5x5�5�5�5�5�56626F6_6t6�6�6�6�6�6	7%7>7R7g7y7�7�7�7�7�7�788'8<8T8�8�8�8�8�8�8�8�89"979K9a9u9�9�9�9�9�9�9	::-:>:P:h:�:�:�:�:�: ;;L;^;p;�;�;�;�;�;<<<4<=<R<g<o<�<�<�<�<�<=*=R=i=�=�=�=�=�=
>>:>Q>p>�>�>�>�>�>??<?Q?l?�?�?�?�?�?   @  h  0080O0n0�0�0�0�0�0�011,1A1U1j11�1�1�1�1�122.272L2a2i2~2�2�2�2�2 3#3F3^3w3�3�3�3�3�34(4<4X4m4�4�4�4�4�45!565Q5h5�5�5�5�5�56646S6l6�6�6�6�6�6�6�67#777L7a7y7�7�7�7�7�7�788(8=8F8Z8r8~8�8�8�8
9)9A9Z9r9�9�9�9�9�9:$:C:X:s:�:�:�:�:�:;$;?;V;u;�;�;�;�;�;<"<A<Z<n<�<�<�<�<�<�<�<=(===R=j=�=�=�=�=�=�=�=>>,>4>I>a>m>�>�>�>�>?/?H?k?�?�?�?�?�?�?   P  d  
0&080M0a0z0�0�0�0�0�01$1@1U1p1�1�1�1�1�1	2"262K2`2t2�2�2�2�2�2�2�23#3;3q3�3�3�3�3�3�3�3�3	4424H4\4u4�4�4�4�4�4�455%5C5R5w5�5�5�56e6w6�6�6�6�6�6�6�67M7`7r7�7�7�7�7�78'898A8S8e8n8�8�8�8�8�899a9s9�9�9�9�9�9�9::0:B:T:n:�:�:�:�:�:�:1;I;[;};�;�;�;�;�;<<(<=<N<l<{<�<�<�<�<�< =5=J=_=h=|=�=�=�=�=>>*>F>r>�>�>�>�>�>�>??,?@?T?m?�?�?�?�?�?�? `  D  	0$0\0n0�0�0�0�0�0�0�0�01121F1_1q1�1�1�1�1�1�1�12!292^2o2�2�2�2�2�2�23303W3i3{3�3�3�3�3�3�3�4�4�4�4�455,5A5V5g5y5�5�5�5I6[6m6u6�6�6�6�6�677&787J7t7�7�7�7�7�7�7!838g8�8�8�8
9959[9�9�9�9::-:B:K:a:u:�:�:�:�:�:�:;';8;J;_;w;�;�;�;�;�;�;<&<S<f<u<�<�<�<�<
=='=@=X=p=�=�=�=�=�=�=�=>)>;>D>Z>n>�>�>R?�?�?�?�?   p  �   0)0L0�0�0�0�0,1>1R1�1�1�1�1U2v2�23V3h3~3�3�3�3�3.4@4R4z4�4�4�4�455_5t5�5�5�5646B6Z6�6�6�67,7@7U7g7�7�7�7�78%898K8�8�8�8�8	9939;9j99�9�9�9�9::::�:;B;`;s;�;$<<<k<}<�<�<�<�<�<e=�=�=�=>,>I>? �  |   ,3K3B4�67J7}7�7�7�7�788<8�8�8�8�8�8�899(9?9T9l9�9�9�9�9�9:#:7:I:i:�:�:�:�:�:;a;�; <�<�<e=z=�= >�>�>9?I?�?�?   �  |   00�0�0�0\2f2�2 44�4�4�466?677)7<7�7�79|9:p:�:�:�:�:�:;4;S;w;�;:<c<�<�<�<=B=e=�=>1>d>�>�>�>?#?^?�?�?�?   �  �   D0�0�0�0111C1~1�1�12d2�2�2�2)3_3�3�3�3�3"4E4�4�4"5M5�5�5�5V6k66�6%797p7�78&8B8W8p8�:�:+;@;U;];s;�;�;�;�;�;<.<C<�<�<=9=�=�=�=�=�=>!>6>J>f>}>�>�>�>�>�>R?~?�?�? �  �   ?0k0 2�2�2�2�2
3�3�3�4i5~5�5�5�5�5�5�556J6_6s6�6�6�6�677�7�7E8e9�;<d<�<T=_=�=�=�=�=>j>~>�>�>�>�>?)?>?S?g?|?�?�?�?�?�?   �  �   0&0t0�0�0�0�0I1�1�1�1�12p2�2�2383�3�3�3�3:4V4�4�4�45.5�5�5�5{6�6�6�6777L7U7i7~7�7�7�78808X8j8�8�8�8�8�8H9]9r9�9�9&:;:�:�:;e;�;�;<:<�<�<�<=�=@>T>h>q>�>�>�>�>
??3?H?]?t?�?�?   �  �   *12"262>2S2g2p2�2�2�2 33)3W3�3�3�3�3�3�3�34Z4n4�4�4�4�4�4�45'5�5�5A6W6�7�7�7�7b89\9g9�97:?:I:y:�:�:�:;C;e;�;E=@>�>F?�?�?   �  �   0j0�0Z1e1J2_2|2�2�2�2�23 353�3�3�3�374L4c4�4�4(5C5X5a5u5�5�5�5�56'6N6�6�6�6�6�67'7<7P7e788+838H8]8f8z8�8�8�89'9�9�:/;=;R;f;�;�;�;�;�;�;d=w=3>A>W>l>�>�>�>�>   �  H   	00d0o0�0�0�01�1�1 22�2�4�4�56U7�7#8`8�839:9l9�9�9n;y;m<V?f?   ,   �1�1�1�1�57(7�7&969�9�9�:;<(<�<=      717579�9:!:5:B;a;u;�;     T   Y021�2�2�2*3A3L3y3�3�3�3�3�3�3�34f4s4�425V6h6787N7d7r7�7�7�78�8�8:(:== 0 X   u0|0�0�0�0�0�01#171�1�1�2�2�2�2*3�5V6e6�7&888D95;<;H;�;�;�;�;�;<h<�<�<�=>>�? @ �   �1�148Q8]8g8�8�8�89909B9�9�9�9�9�9::A:R:t:�:�:�:�:�:�:;;1;B;d;�;�;�;�;�;< <0<T<t<�<�<�<�<�<�<= =/=?=P=�=�=�=�=�=>$>D>d>�>�>�>�>�>?4?d?�?�?�?�? P    00D0a0t0�0�0�0�01!111D1d1�1�1�1�12$2D2d2�2�2�2�23353'4X4j44�4�4�4D5o5�5�5�56$6D6d6�6�6�6�67!747d7�7�7�7�7�788-8;8J8\8�8�8�8�8�89$9Q9a9q9�9�9�9�9�9�9�9::,:T:t:�:�:�:�:;4;T;t;�;�;�;�;<)<E<]<w<�<�<�<�<=4=T=t=�=�=�=�=�=�=>">1>A>S>t>�>�>�>�>�>?"?7?Q?b?�?�?�?�?�?�?   ` �   40T0t0�0�0�0�011$1D1d1�1�1�1�12$2D2d2�2�2�2�23$3D3d3�3�3�3�34$4L4t4�4�4�45$5D5d5�5�5�5�56$6D6d6�6�6�6�67$7D7d7�7�7�7�78!848T8t8�8�8�8�8�89949T9v9�9�9�9�9	:*:d:�:�:�;�;�;�;�; <5<�<�<�<�<=$=T=t=�=�=�=>4>F>t>�>�>\?�?�?�?�? p �   70w0E1J1U1x1�1�1�1�12A2t2�2�213d3�3�3�3*4V4k4�4�45K5�5�5�5 6P6�6�6�6�6�6767M7w7�7�7�7818P8l8�8�8�89/9k9�9�9�9�9:G:q:�:�:�:;;g;�;�;�;�;*<�<�<�<�<U=�=�=K>�>�>�>(?k?�?�?   � �   	0#0l0�0�0161Q1�1�1�12d2�2D3�3�3$4f4x4�4�4N5m5�5!6]6�6�6�6+7G7_7v7�7�7�7*8J8�849y9�9 :c:�: ;S;�;<s<�<=s=�=3>�>�>S?�? � �   0s0�0#1�1�1I2�2�2Y3�3 404j4�4�4�4 5T5~5�5616k6s6�6�67J7�7�78~8�8�8>9t9�9�9:A:t:�:�:$;a;�;�;�;<4<a<=
==+=H=R=�=�=.> ?�?�?�?�?�?�?�?�?�?�? � �   &0�0014181<1@1D1H1L1P1�12"2D2o2�2�2�2�23!3A3d3�3�3�3444d4�4�4545a5�5�5T6t6�6�6�6747d7�7�7�7868H8Z8x8�8�8�8�8�89 919E9c9|9�9�9�9�9�9�9$:t:�:�:�:;T;�;�;�;$<<<�<�<�<$=Q=�=�=T>�>�>�>�>%?�?�?�? � �   0"0�041�1�1�1�1�12242�2�2�2363J3Z3�3�3�3C4�45i5�5�5�5$6Q6�637c7�7�7�7�718F8Z8o8�8�89A9x9}9�9�9�9�9:D:A;;�;�;�;�;<%<`<�<�<�<�<�<*=N=g=�=�=�=>">I>�>�>�>�>�>�>?/?O?m?�?�?�? � �   0@0v0�01�1�1�12C2m2�2�2�2"3T3�3�3�3�34494G4g4{4�4�4�4�4�45545O5a5t5�5�5�5�5�5�7~8�89T9�9):�:�:$;E;�;�;d<�<8=Y=>>F>Y>k>|>�>�>�>	?&?Y?�?�?�? � �    00O0a0s0�0�0�0�0-1;1K1�2�2�23[3w3�3�3�34A4l4�4�4�4C5U5�5�596U6�6�697\7x7�7�7�7�78}8�89l9�9�9:4:T:t:�:�:�:�:;4;d;;�;�;�;�;!<4<d<�<�<�<=!=D=t=�=�=�=>4>a>�>�>�>?$?D?d?�?�?�?�? � �   0$0D0a0t0�0�0�0�0^1~1�1272�2�23�3�3�3H4j4�45565�5�5�5c6�6�6�67T7�78D8�8�89�9�9�9^:~:�:;|;�;<'<�<�<='=�=�=c>�>�>.?N?c?�?�? � �   0a0w0�0<1�1�1�12!242d2�2�2�2�2343q3�3�3�3�3444g4�4�4�45>5W5k5�5�5�5616T6q6�6�6N7S7X7]77�7�7�78$8D8d8�8�8�8949T9t9�9�9�9�9�9:R:�:�:�:";P;~;�;�;�;<$<T<�<�<�<�<=D=d=�=�=�=>D>d>�>�>�>�>?$?D?V?q?�?�?�?�?�?     �   0$0D0�0�0�0�01$1D1d1�1�1�1�1�1�1242T2t2�2�2�23$3D3a3t3�3�3�34444�4�4�4�4545T5t5�5�5�5�5646t6�6�6#7s7�7�7!8D8t8�8�8�89$9A9Q9d9�9�9�9�9:9:M:�:�:�:;4;T;t;�;�;�;�;$<B<V<f<�<�<�<�<=4=`=t=�=�=�=�=>:>m>{>�>�>�>�>�>?$?>?R?b?�?�?�?�?    �   0,0U0�0�0�0�0�0�0%1S1i1w1�1�1�122T2}2�2�2�2343_3�3�3�3�34$4A4T4t4�4�4�45$5D5d5�5�5�5�56$6D6a6q6�6�6�6�67717T7i7{7�7�7�7�7�8�8959u9�9�95:�:�:�:;E;�;�;<M<�<�<=R=�=�=>E>�>�>?R?�?�?�?     �   20e0�0�051u1�1�182S2�2�2�2�23U3�3�34e4�4�4A5i5�5�5�5�5�56B6j6�6�6�67X77�7�7"8e8�8�8�89R9�9�9�98:v:;2;G;d;�;�;�;�;<!<1<D<a<q<�<�<�<�<�<=4=T=t=�=�=�=�=>D>d>�>�>�>�>?$?D?�?�?�?�?�? 0 �   0!0?0a00�0�0�0111T1t1�1�1�1�12$2A2T2t2�2�2�23$3D3�3�3�3�3!4A4a4�4�4$5t5�5�5�5646T6t6�6�6�6�6$7D7t7�7�7�7848a8�8�8�8919T9�9�9�9:1:Q:q:�:�:�:�:;1;Q;q;�;�;�;�;<1<Q<t<�<�<�<=$=D=a=�=�=�=�=>>A>a>�>�>�>�>?$?D?t?�?�?�?�? @ �   040k0�01R1�1�1�12$2T2�2�2�2�2343a3�3�3�3444~4�4�45$5D5d5�5�5�56!6A6d6�6�6�6747d7�7�7�7�7818D8a8�8�8�8$9�9�9�9�9:4:d:�:�:�:;1;Q;q;�;�;<$<D<t<�<�<�<$=d=�=�=>A>a>�>�>�>?$?2?7?T?}?�?�?   P �   *0T0t0�0�01W1�1W2�2�2�2�2343]3�3�3�3$4A4d4�4�4�4�5�5�56$6T6�6�6�6�6747R7s7�7�7�7848Q8t8�8�8919T9�9�9�9�9!:4:T:�:�:;1;T;t;�;�;�;<a<~<�<�<�<=2=[=l=�=�=�=�=>&>N>b>�>�>�>?%?[?n?�?�?�?�?�?   ` t   �0�011T1\1�1�1�3�6�6�67@7P7�7�7�7�9�9�9�9�9�9:8:�:;�;�;<'<�<�<D=�=�=>!>1>M>q>�>�>??9?U?v?�?�?�?�?   p   0M0a0q0�0�0�0�0
1'1X1�1�1�1�1�1$2w4�41585w5�5�5
66D6M6Z6t6�6�6�6�6�6�6�6�6757G7b7x7�7�7�7�7�7�78)8;8M8_8h8�8�8�8�8�899(919O9p9�9�9�9�9�9::':9:K:]:o:x:�:�:�:�:�:;&;8;A;_;�;�;�;�;�;�;�;<4<_<�<�<�<�<�<�<�<�<=&=D=V=r=�=�=�=�=�=�=>&>B>T>f>o>�>�>�>�>�>?'?9?V?l?�?�?�?   � �   0r0z0�0�0�0�0�0�01
11o1�1�1�1�1e2w2�2�2�2�2343T3h3z3�3�3�344�4�4�4A5�5�5�5�5�56$6D6a6t6�6�6�6�67,7�7�8�8�8�8�8�8�8�8�8�89I9�9u:�;�;<�<===%=,=3=:=A=H=O=V=]=d=k=r=y=�=??4?A?G?s?z?�?�?�?�? � �   0(0,0004080<0X0f0�0�0)1�1�1�1�1�12h2�2�2�2�2
3t3�3�3�3�3!4d4�4�4�4�4�45505\5�5�5�5�5�5+6:6r6�6�6�6�6�6�637L7y7�7�7�7,838 � (   �2�<=-=e=�=�=5>u>�>�>"?U?�?�?   � p   0E0�0�0121b1�1�1�152u2�23U3�3�34e4�4%5u5�5�5E6(8G8�:H;L;P;T;X;;<I<h<v<==5===�=>0>>>w>�>�?�?�?�?   � �   @0N0c0q0Q1d1�1�1�1�12D2c2v2�2�2�23A3T3�3�3�3�34$4T4�4�4�4�4$5d5�5�5�5�56$6D6t6�6�6�6a7t7�7�788(:::M:p:>;V;�<=$=T=�=�=�=�=�=>#>D>d>�>�>�>??$?Q?t?�?�?�?�?   � d   0D0(1\1�1�1+2�233�3�3�324�4�45$5U5�5�5G6X6*:�:�:�;0<�<�<�<�<====�=�=�?�?�?�?�?�?�?�?   �   0+0�0�0�0�0�0�0�01}1�1�1�1�1�12)222K2[2{2�2�2�233#3(3h3�3"4+4�5�5�5�5�56)636P6p6�6�6�6�6?7�7�7�7�7�7�7�7�7888�8A9I9^9i9�9r;7<p<�<�<�<�<�<�<�<�<�<�<�<======"=&=?=z=�=�=�=�=�=�=�=>3>Q>X>\>`>d>h>l>p>t>�>�>�>�>�>6?A?\?c?h?l?p?�?�?�?�?�?�?   � �    00000Z0`0d0h0l0 11f1�1�1�122I244�4�4�45 585x5�5�5�566.6�6J7b7g7�9�9*:�:�:�:�:.;�;�;�;�;O<m<�<+=M>p>{>�>�>'?�?     �   80�1]3�4�5�5�6�6�6�6$7<7D7J7�7�7�7�7�78h8�89J9c9�9:
::2:N:�:�:@;F;f;�;�;�;J<<�<�<�<�<�<�<�<=!=(=,=0=4=8=<=@=D=�=�=�=�=�=>>,>3>8><>@>a>�>�>�>�>�>�>�>�>�>�>*?0?4?8?<?�?�?  �   0.0W0\0s0�0�0�0P1b1�1�1�1�1�1�1�1222K2{23�3�3c445�5�556A6�6�637?7�7�788D8h8J9�:�;�;�;�;<<3<;<g<p<|<�<�<�<=
==S=\=h=>">E>	??+?=?[?�?�?   t   �0�01^1�1�1�2�2�2�2333*363B3N3Y34�4�4!5t5z5�5�5�566o6�6?7@8�8�:;K;�;�;�;d<�<�<�<>�>�>�>�>??u?�?   0 �   �01�1�344:5w5�577L7Y7c7q7z7�7�7�7�7�7�78'8^8�8�8939{9�9:{:�:�:�:�:�:�:�:;#;,;2;;;@;O;v;�;�;�;�;�;�;�;�;<<><D<O<[<p<w<�<�<�<�<�<�<�<�<�<�< ====%=/=6=N=]=d=q=�=�=�=>>?>E>a>y>�>?<?F?~?�?�?�?�?�?�?   @ �   
00%030>0E0`0e0m0s0z0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0111(1-181=1J1X1^1k1�1�1�1�12/2B2�2�2�2�2�2�2�2�2�2�2�2�2�2�2333$3)3/393B3M3Y3^3n3s3y33�3�3�4@5�798q8�=�>   P �   *0x0�0�0�0�0�0A2^2c2q2y2�2�2�2�2�2�2�2�2�2�2�2�2�23-3;3A3d3k3�3�3�3�3�3�3s4�4�4�4�6�6�677+747A7L7^7q7|7�7�7�7�7�7�7�7�7�7�7�7�7�78	888#8,898?8Y8j8p8�8�8�<�<�<�<!=f=9?D?L?a?~?�?   ` X   �0�0�0�0;1_1l11G2m3f4�4K6�7�:	;;=>T>_>�>�>�>�>??)?5?E?L?[?g?t?�?�?�?�?�?�? p t   00?0H0l0�0`1v1�1�12
2<2�2�2�2�23&3g3�3�3�34%4C4e4�5�56]6�6v7�7�8�89�:v;?<p<�<�<�<�=�=�=_>�>�>�>�>~?�?   � 8   �0A1�253B3b3|3�3�3�4S5�6�617;7S7|7�7�79�9�9�9   � d   �0;;5;>;k;�;�;�;�;�;<%<8<C<H<X<b<i<t<}<�<�<�<�<�<�<�<1=>=h=m=x=}=�='>4><>K>�>�>�>�>�>?? � �   �0�0�0�0�0�0W1]1s1~1�1�1�1�1�1;2N2�2�2�2�2�2�23�3�3�3�3y4�4�4�4�4�4�4�4�465>5K5�5�56!6<6H6T6`6�6�6�6�6�6�6�6�6�6777%717:7C7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7=8�8�89949=9D9M9�9�9�9�9::/:A:e:�:�:�;�;�<�<==S=�=�=�=>�>!?1?=?O?_?k? � <   i0�0x1�182~2�2�2�23035:y;�;�;�<�<�<�<1>L>�>A?K?m?   � �   ;0<1L1]1e1u1�1�1�1�12$233I4S4k4r4|4�4�4�4�4a5�5@6�6�6�6�6	7^7�7�748:8�8�8�8�8999e9�9�9:	::H:V:�:�:�:�:�:�:�:;s;|;�; � h   �12=2O2a2�2�3�3�3�3M4_4q4�4�4�4�4�4�6?7P7v9�9�9�9�9�9::�:�:%;I;�;�;k=�=c>l>�>�>?E?�?�?�?�?   �    0@0O0�5 � x   �6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�677777777#7'7+7/737�7I9�9�9�9:7:Y:d:�:�:�:�:�:; ;%;�;�;�<�>�>_?     h   ~1�3�3�3�3�4�4�4�4�4�4l5�5�5U6o6x6�6�6�6�6�6 77v7�759�9�9�:�:1;>;< <�<�</=^=9>F>_>}>�>�>�?�?    �    000#0A0K0T0_0t0{0�0�0�0W1�1�12!2F2�2�2�2�2"333n3�3�3�34,454u4�4�4�45P5X5�5n69k:�:�:�:�:%;.<�<�<4=�=�?�?�?�?�?�?     x   (0b0p0v0�0�0�0�0�0�0�0�0�0�0�0�011V1s1�1�1�1�1�2T3r3�3�34&4q7a8�9:?:"<>">&>*>.>2>6>:>_>z>�>�>�>�>�>�>|?�?   0 @   0 1E2�3u6�6`7s7�7�7�7�78&8	;+;c;�;�;�;�;�;<�<�=�>�?   @ @   �0�0n1P2�2�2�3�3�3G4^45�5�5�6�7-838�8�8�8�9�9�9_:/=F=   P D   �0�0�0�0�0�0�0�0�0�0�0�0�0�1�1�1�1Y2}2�<4>:>?>E>L>^>r>}>�?�? ` l   �0�0_1f1�1�1<23�34!666R6r6�6�6�6�67E7b7�7�7�7�78?8b8�8�8�8�899'939?9I9U9b9j9t9�9�9�9�9�9�9�9   p �  `1d1h1l1p1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8�8�8�:�:�:�:�:�:�:�:�:�:�;�;�;�;�;�;�;�;�;�;<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=�=�=�=�=�=l>p>8?<?@?D?H?�?�?   � d   H0L0P0T0X0\0`0d0t0x0|081<1@1D1H1L1P1T1l1p1t1@:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�;�;�;�;�;�;   � �   �9�9�9�9�9�9�9 :::: :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�< � x  �2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3d6h67777 7(7@7D7\7l7p7�7�7�7�7�7�7�7�7�7�7�78888$8<8L8P8T8\8t8�8�8�8�8�8�8�8�8�8�8�8�8�89$9(909H9X9\9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9::,:<:@:P:T:d:h:l:p:x:�:�:�:�:�:�:�:�:�:�: ;;;$;4;8;H;L;P;T;\;t;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<(<,<<<@<D<L<d<t<x<�<�<�<�<�<�<�<�<�<�<�<�< ===$=(=,=0=8=P=`=d=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=>>$>(>8><>@>D>L>d>t>x>�>�>�>�>�>�>�>�>�>�>�>�>?? ?0?4?8?@?X?h?l?|?�?�?�?�?�?�?�?�?�?�?�?   � �   000$04080H0L0P0X0p0�0�0�0�0�0�0�0�0�0�0�0�0�01$1(181<1D1\1l1p1�1�1�1�1�1�1�1�1�1�1�1 22222$2<2L2P2`2d2h2l2t2�2�2�2�2�2�2�2�2�2�2�2333343D3H3X3\3`3h3�3444 4(4<4D4X4h4�4�4�4�4�4�45(5<5L5p5|5�5�5�5�5�5�5 6,646L6T6\6`6d6l6�6�6�6�6�6�6�6�6�6�677747<7D7H7L7T7h7p7�7�7�7�7�7�78 808\8d8�8�8�8�8�8�89(949<9\9�9�9�9�9�9�9�9:0:<:D:d:t:�:�:�:�:�:�:; ;@;H;T;t;|;�;�;�;�;�;�;�;�;�;<(<H<h<�<�<�<�<�<=0=P=l=p=�=�=�=�=�=>(>H>h>�>�>�>�>�>�>�>?8?@?D?\?`?p?�?�?�?�?�?�?�?   � X    00 0(00080<0D0X0t0x0�0�0�0�0�0�0181X1x1�1�1�1�1282T2X2t2x2�2�2�2�23$3<3@3`3 � $   00 080<0@0\0x0�0�0�0�01L1�1�1�102P2�2�2 3 3@3d3�3�3�3�3�3�34 4$4(4,4H4d4|4�4�4�4�4�4�4�4�4�4�4�4�4�455 5$5(5,5054585<5T5X5\5`5d5h5l5�5�5�5�5�5�56 6$6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�607P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�;H=X=h=x=�=�=�=�=�=�=�=�=�=P?T?X?\?`?d?h?l?p?t?   � p  �0�0�0�0�3�3�3�3�3�3�3�3�3�3�3�34444$4,444<4D4L4T4\4�4�4�4�4�455
555555"5&5*5.52565:5>5B5F5J5N5R5V5Z5^5b5f5j5n5r5v5z5~5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�68$8,848<8D8L8T8\8d8l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8D9H9�9�9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                