MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��."��@q��@q��@q$��q��@q��q��@q��q'�@q���q��@q��Aq�@q��q�@q��q��@q��q��@qRich��@q                PE  L ���Q        � !
  D  �      v     `                       `         @                    � S   �� <                             �7  �a                            @� @            ` H                          .text   �C     D                   `.rdata  sg   `  h   H             @  @.data   D:   �     �             @  �.reloc  :C     D   �             @  B                                                                                                                                                                                                                                                                                                                                                                                                U��Ejj j P��M ��]����������U��]�N �������U�졸�V��H�QV�ҡ���U�H�E�IRj�PV�у���^]� ����������U�졸��P�E���   ��VWP�EP�E�P�ҋu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]� ������������V���Xw �N��a�r �N$�N ��^���������������V��N$��a��N �N��r ��^�?w ���������������U���T  ���3ŉE�Wj j�WK ����u_�M�3���� ��]�V������PWǅ����(  �$K ����   ������Qj�K �����   ������RPǅ����$  ��J ���}   ������P������h  Q�� ������h  R�� ���������P�I �@��u�+�$    ��/t��t������H��\uꍴ����V�[� h bV�� ����u.������PW�PJ ���8���W� `^3�_�M�3���� ��]ËM�^3͸   _��� ��]���������3���������������3������������������������������j j j�� �����U���lV��E�P�M�Q���E�   �E�    �� �}� �f  SW�M���K ����B�P�M�Q�ҡ���P���   ���E�Pj�M̍~Q���ҋء���H�A�U�R�Ћ���Q�J�E�PS�ы���B�P�M�Q�҃��E�P�M���K �M�Q�M���O �M��WL ����B�P�M�Q�ҡ���H�A�U�R�Ѓ�h�b�M��dK �M�Q�M���O �M��L �U�j R�%] �����f  ����H�A�U�R�Ћ���Q�Jj j��E�h�bP�эU�R�  ����H�A�U�R�Ѓ�j ���Hw ����Q�J�E�P�ы���B�Pj j��M�h�bQ�ҍE�jP��� ����Q�J���E�P���у� ����   ����B�P�M�Q�ҡ���H�Aj j��U�h�bR�ЍM�Q��� ����B�P�M�Q����� jh(bh�   h�   ����H ��,��t	���K�  �3�WS���N�  h�  ���bv �M��J _[^��]� j j �E�P���E�   �E�    �� �M��J _[^��]� ���U���SVW��j�~W�E�3�P�E�   �]��� jW�M�Q���E�   �]��� jW�U�R���E�   �]��*� jW�E�P���E�   �]�貀 jW�M�Q���E�   �]�蚀 jW�U�R���E�   �]�肀 jW�E�P���E�   �]��j� jW�M�Q���E�   �]��R� j
W�U�R���E�
   �]�蚀 j	�E�	   �]�W�E�P���"� jW�M�Q���E�   �]��
� jW�U�R���E�   �]��� jW�E�P���E�   �]���� jW�M�Q���E�   �]��� _^[��]������������U���   V����� ��u^��]�SWhc�M��'H �E�P�M�Q�~$��] ��P�U�R��L ��P���L �M��H �M��H �M��H 3ۉ^@�_ SW�E��Y �����z  �E�P���=I P�M���G jj�M�Q�M�htaoc�_ ���M��E��QH ����B�P�M�Q�҃�8]�t�E�P�^_ ��_[3�^��]Ë���Q�J�E�P�ы���B�PSj��M�hcQ�ҡ���P�R8���E�P�~j���ҡ���H�A�U�R�Ѓ��M���F �M�j	Q�] ��P�M��xK �M��G hc�M���F h�b�M���F �U�R�E�P�M�Q��l���R�nK ��P�E�P�aK ����l����SG �M��KG �M��CG �M�jQ�XX ����t6�U�R�M���G ����QP�B8j���Ћ���Q�J�E�P���   ����B�P�M�Q�ҡ���H�ASj��U�h�bR�ЍM�Q�� ����B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�JSj��E�hcP�ы���B�P8��0�M�Qj���ҡ���H�A�U�R�Ћ���Q�B4��Sj���Ћ���Q�B0jj���Ћ���Q�B0jj���Ћ���Q�B0Sj���Ћ���Q�B0Sj���Ћ���Q�B0jj���Ћ���Q�B4Sj
���Ћ���Q�B0jj	���Ћ���Q�B0jj���Ћ���Q�B0Sj���Ћ���Q�J�E�P�ы���BSj��P�M�hcQ�ҡ���P�R8���E�Pj���ҡ���H�A�U�R�Ћ���Q�B0��Sj���ЋM�W�c �M��\ �M��E �M��E �M�Q�N$��E P�M��yD �M�jj�U�Rhtaoc�D\ ���M��E���D ����H�A�U�R�Ѓ�8]�t�M�Q��[ ��_[3�^��]ËM�j�~W��^ �M��\ ����E�   �]�B�P�M�Q�҃�SS�E�Pj�M�Q�������P�U�R���v ����H�A�U�R�Ћ���Q�J�E�P�ы���E�   �]�B�P�M�Q�҃�SS�E�Pj�M�Q������P�U�R���Sv ����H�A�U�R�Ћ���Q�J�E�P�у��E�   �]�h�������B���   h  �Sjh���h  �Sj����P�E�P���
q ���S�E�   �]�Q���   Sj����P�M�Q���ݽ ���S�E�   �]�B���   Sj����P�E�P��谽 ���S�E�   �]�Q���   Sj����P�M�Q��能 ���S�E�   �]�B���   Sj����P�E�P���V� ����E�   �]�S�Q���   Sj����P�M�Q���)� ���h���h  �Sjh���h  ��E�
   �]�B���   Sj
����P�E�P����o ���S�E�	   �]�Q���   Sj	����P�M�Q��蹼 ���S�E�   �]�B���   Sj����P�E�P��茼 ���S�E�   �]�Q���   Sj����P�M�Q���_� ����E�   �]�B�M̋PQ�҃�SS�E�Pj�M�Q���-���P�U�R���t ����H�A�U�R�Ћ���Q�J�E�P�ы����S�E�   �]�B���   Sj����P�E�P���λ h�  ����l �M�Q�iX ��_[�   ^��]�����������U���0V��~@ t~W�+X �E��E�P�N$�A P�M��s@ jj�M�Q�M�htaoc�>X �MЋ���@ ����B�P�M�Q�҃���_t���3����M���V�^ �M��X �E�P��W ��^��]���������������U����   SV��3�W�]��F@   ������E����   ����   H��  ����H�A�U�R�Ћ���Q�JSj��E�h�bP�эU�R��� ����H�A�U�R����� jh(bh  h�   ����= ��,;�t���E�  ��VW���I�  _^�C[��]� ��3�VW���/�  _^�   [��]� �MQ�U�R���E�   �]��xt 9]��  h�  ���k _^�   [��]� �P� jh(bh�   j$���[= ��;�t�@   ��X�X�X�X�3���VW���U  ����H�A�U�R�Ћ���Q�JSj��E�hTcP�эU�R�� ����H�A�U�R�Ћ���Q�J�E�P�ы���B���   �� �M�Qj��8���R���Ћ���Q�J���E�P�ы���B�P�M�QW�ҡ���H�A��8���R�Ћ���Q�J�E�P�ы���B���   ��Sj���҅�tR����H�A�U�R�Ћ���Q�JSj��E�hcP�ы���B�Px���M�Q�M��E�   ���E��u�]�E�t����H�A�U�R�Ѓ�8]�/  ��������   ����Q�Bdj�M��Ћ���Qh(b�p���   h�   V�Ћ���Q��j���BhVW�M���j<��H���SQ��� ����H���RǅH���<   ��L�����P���ǅT���Lc��X�����`���ǅd���   ��h����@a��uwSh4c�M��=����E�P��� ����Q�J�E�P�у��I����B�P�M�Q�ҡ���H�ASj��U�h cR�ЍM�Q�y� ����B�P�M�Q�҃�����H�A�U�R�Ѓ�_^�   [��]� ��U��V��N$��a�\< �N�d` ����d �Et	V�; ����^]� �������U��M�U�A�
�E��B�I0���B�IH����A �
�A�A8�J���AP�J���X�A(�
�A�A@�J���AX�J���X�A�J�B �I0���B(�IH���X�A8�J �A �J���AP�J(���X �A@�J �A(�J���AX�J(���X(�A�J0�A0�J8���AH�J@���X0�A8�J8�A �J0���AP�J@���X8�A@�J8�A(�J0���AX�J@���X@�A�JH�BP�I0���BX�IH���XH�BP�I8�BH�I ���AP�JX���XP�A@�JP�BH�I(���AX�JX���XX]���U�졸��H�U�I(��VWR�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]���U���$�ESVW3ۍM�Q�M��]܉]�E�]��]��' �}S�U�R�E�P��� �M����	 ;�th������   �JX�E�P�ы���;�tJ������   �PT���ҋ���Q|�M�RQPV�ҋ�����   ��U�R�Ѓ�_��^[��]� ������   �
�E�P�у�_^3�[��]� ������������U���$�EVW3��M�Q�M��}܉}�E�}��}��H �MW�U�R�E�P�� �M����= ;�tZ������   �JH�E�P�ы���u���B�HV�ы���B�HVW�ы�����   ��M�Q�҃�_��^��]� ����H�u�QV�ҡ���H�QWj�hcV�ҡ�����   ��U�R�Ѓ�_��^��]� ��������U���$�EVW3��M�Q�M��}܉}�E�}��}��X �MW�U�R�E�P�� �M����M ;�t8������   �J8�E�P�ы�������   ��M�Q�҃�_��^��]� ������   ��U�R�Ѓ�_3�^��]� �U���$�ESV3��u��M�Q�M��u܉u�E�u��u�� �MV�U�R�E�P�4 ��t ������   �J�E�P�у���t��2ۍM�� ^��[t7������   �P<�M�Q���]������   ��U�R���E����]� ������   �
�E�P���E����]� ���������U���$�EVW3��M�Q�M��}܉}�E�}��}��� �MW�U�R�E�P�g �M����� ;�t[������   �J@�E�P�ыu��H��P�N�H�V�P�@�N����V���   �
�F�E�P�у�_��^��]� �����u����   �V��^�M�Q�҃�_��^��]� U���$�EVW3��M�Q�M��}܉}�E�}��}�� �MW�U�R�E�P� �M���� ;�tD������   �JL�E�P�ыu��P����5 ������   ��M�Q�҃�_��^��]� �uW���*5 ������   ��U�R�Ѓ�_��^��]� ����������U��Q����P�BdVWj�M�Ћ���Qh�c�p���   h�  V�Ћ����j�E��QVP�Bh�M��N3���~S�]�I �M��R���A G;�|�[�E�P�2 ����Q�J�EP�у�_^��]� �����U�������H�AV�U�WR�Ћ���Q�Jj j��E�h�cP�ы���B�Pd��j�M��ҍp����H���   h�ch�  V�ҋ����j�E��QVP�Bh�M���N3���~S�]���M��R����@ G;�|�[�E�P�B1 ����Q�J�E�P�у�_^��]� �����U��Q�ESVW���   3�3�3�3ۉM���|!�@|�O���A�	�d$ p��Iu��E�M�;�}�@|��_�^�[��]� �������U�졸��H�Q��   V�uV�ҡ���H�Qj j�h�dV�ҋE����
�  �$��. j h�d�M�������E�P���m  ����Q�J�E�P����  j h�d��`���������`���R���Wm  ��`����  j hxd�M��}����M�Q���2m  ����B�P�M�Q���p  j htd�M��L����E�P���m  ����Q�J�E�P���?  j hpd�M������U�R����l  �U��  j hhd�M�������M�Q���l  ����B�P�M�Q����   j hdd�M�������E�P���}l  ����Q�J�E�P���   j h\d�M������U�R���Ll  �U��   j hTd�M��u����M�Q���*l  ����B�P�M�Q���kj hLd��p����D�����p���P����k  ����Q�J��p���P���4j hDd��P���������P���R���k  ��P�������H�AR�Ѓ�����Q�J�E�P�ы���B�Pj j��M�h@dQ�ҡ���P�B<�����Ћ���Q�RLj�j��M�QP���ҡ���H�A�U�R�Ѓ���^��]� �I H, y, �, �, - (- Y- �- �- �- . ����S�   V3�W���7�G�w�w�w�w�G(�w�w�w,�w$�w �G@�w0�w4�wD�w<�w8�GX�wH�wL�w\�wT�wP�Gp�w`�wd�wt�wl�wh���   �wx�w|���   ���   ���   �_���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   97t	W��, ���7�w�w�w�w93t	S��, ���G0�3�s�s�s�s90t	P�, ���GH�w0�w4�wD�w<�w890t	P�, ���G`�wH�wL�w\�wT�wP90t	P�, ���Gx�w`�wd�wt�wl�wh90t	P�b, �����   �wx�w|���   ���   ���   90t	P�7, �����   ���   ���   ���   ���   ���   90t	P�, �����   ���   ���   ���   ���   ���   ��_^[����������SVW���� ���   3�93t	S�+ ���3�s�s�s�s9��   ���   t	S�+ ���3�s�s�s�s9wx�_xt	S�p+ ���3�s�s�s�s9w`�_`t	S�Q+ ���3�s�s�s�s9wH�_Ht	S�2+ ���3�s�s�s�s9w0�_0t	S�+ ���3�s�s�s�s9w�_t	S��* ���3�s�s�s�s97t	W��* ���7�w�w�w�w_^[�����U���  ���SVW���H�A�U�R�}��Ћ���Q�Jj j��E�h�dP�ы���B�P�M�Q�ҡ���H�Aj j��U�h�dR�Ћ���Q�E�R(P�M�Q�ҋ���H�A�U�R�Ћ���Q�J�E�PV�ы���B�P�M�Q�ҡ���H�A�UЃ�@R�Ћ���Q�R�E�P�M�Q�ҡ���P���B<�M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ]����Q�B��S����V�Ћ���QV�E��JP�у����P����u�~ �E�    ��  3�����B�P�M�Q�ҡ���H�Aj j��U�h�cR�Ћ���Q�J�E�P�ы���B�Pj j��M�h�dQ�ҡ���H�A��x���R�Ћ���Q�Jj j���x���h�dP�ы���B�P��8���Q�ҡ���H�A��@j j���8���h�dR�ЋF����D8�Q�J$��j0j jj ���������$P�ы��������؋BQ�P�ҡ���H�A�����RS�Ћ���Q�J������P�ыF����D8�B�P$��,j0j jj ���������$Q�ҋء���H�A��(���R�Ћ���Q�J��(���PS�ы���B�P������Q�ҋF�8����H�A$��,j0j jj ��������$R�Ћ���Q�J�؍�H���P�ы���B�P��H���QS�ҡ���H�A�����R�Ћ���Q�J�E�P�ы���B�@�M�Q��8���R�Ћ���Q�B<��8�M��Ћ���Q�RLj�j���H���QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j���x���QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P���B<�M��Ћ���Q�RLj�j���(���QP�M��ҡ���H�A��h���R�Ћ���Q�R��h���P�M�Q�ҡ���P�B<����h����Ћ���Q�RLj�j��M�QP��h����ҡ���H�A��X���R�Ћ���Q�R��X���P��h���Q�ҡ���P�B<����X����Ћ���Q�RLj�j������QP��X����ҡ���H�A�U�R�Ћ���Q�R�E�P��X���Q�ҡ���P�B<���M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A��X���R�Ћ���Q�J��h���P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P��H���Q�ҡ���H�A��(���R�Ћ���Q������JP�ы���B�P��8���Q�ҡ���H�A��x���R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҋE����Q��<P�B����S�Ћ���Q�J�E�SP�ыM̃�������E�@���E�;F�u����}̋]����B�P��x���Q�ҡ���H�Aj j���x���h�dR�Ћ���Q�J�E�P�ы���B�Pj j��M�h�dQ�ҡ���H�U�I(R�����P�ы�����B�P�M�Q�ҡ���H�A�U�RV�Ћ���Q�J�����P�ы���B�P�M���@Q�ҡ���H�I�U�R�E�P�ы���B�P<���M��ҋ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j���x���QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҡ���H�A��x���R�Ћ����S����Q�BV�Ћ���Q�J�E�VP�у�������S���;�������B�P�M�Q�҃�_^[��]� �������������U���  ���SVW���H�A�U�R�}��Ћ���Q�Jj j��E�h�dP�ы���B�P�M�Q�ҡ���H�Aj j��U�h�dR�Ћu�F,����Q�J(P�E�P�ы���؋B�P�M�Q�ҡ���H�A�U�RS�Ћ���Q�J�E�P�ы���B�P�M���@Q�ҡ���H�I�U�R�E�P�ы�����B�P<�M��ҋ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�ЋM����B��Q�H����S�ы���BS�P�M�Q�҃�������3ۉ]9]��  ����H�A��(���R�Ћ���Q�Jj j���(���h�cP�ы���B�P������Q�ҡ���H�Aj j�������h�dR�Ћ���Q�J������P�ы���B�Pj j�������h�dQ�ҡ���H�A��h���R�Ћ���Q�J��@j j���h���h�dP�ыF�����j0j �<[�j���D8�B�P$j ���������$Q�҉E�����H�A������R�Ћ���Q�M��R������PQ�ҡ���H�A������R����F�d8����Q�J$��,j0j jj ���������$P�ы���E��B�P������Q�ҡ���H�E��I������RP�ы���B�P������Q�ҋF�8����H�A$��,j0j jj ���������$R�Ћ���Q�J�E���H���P�ы���B�U��@��H���QR�Ћ���Q�J������P�ы���B�P��x���Q�ҡ���H�I��x���R��h���P�ы���B�P<��8��x����ҋ���Q�RLj�j���H���QP��x����ҡ���H�A������R�Ћ���Q�R������P��x���Q�ҡ���P�B<���������Ћ���Q�RLj�j�������QP�������ҡ���H�A������R�Ћ���Q�������RP������Q�ҡ���P�B<���������Ћ���Q�RLj�j�������QP�������ҡ���H�A������R�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j�������QP�������ҡ���H�A������R�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j�������QP�������ҡ���H�A�U�R�Ћ���Q�R�E�P������Q�ҡ���P�B<���M��Ћ���Q�RLj�j���(���QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A������R�Ћ���Q�J������P�ы���B�P������Q�ҡ���H�A������R�Ћ���Q�J��x���P�ы���B�P��H���Q�ҡ���H�A������R�Ћ���Q�J������P�ы���B�P��h���Q�ҡ���H�A������R�Ћ���Q�J������P�ы���B�P��(���Q�ҋE����Q��<P���ĉE�P�B�Ћ���Q�E��RP�M�Q�ҋM�����������H�A��x���R�Ћ���Q�Jj j���x���h�cP�ы���B�P������Q�ҡ���Hj �Aj�������h�dR�Ћ���Q�J������P�ы���B�Pj j�������h�dQ�ҡ���H�A�����R�Ћ���Q�J��@j j������h�dP�ыV�D:(��j0j �D:����H�A$jj ����X����$R�Ћ���Q�J�E�������P�ы���B�U��@������QR�Ћ���Q�J��X���P����V�d: �D:����H��,�A$j0j jj ��������$R�Ћ���Q�J�E���8���P�ы���B�U��@��8���QR�Ћ���Q�J�����P�ыV����D:�H�A$��,j0j j�|:j ����8����$R�Ћ���Q�J��������P�ы���B�P������QW�ҡ���H�A��8���R�Ћ���Q�J��h���P�ы���B�@��h���Q�����R�Ћ���Q�B<��8��h����Ћ���Q�RLj�j�������QP��h����ҡ���H�A��(���R�Ћ���Q�R��(���P��h���Q�ҡ���P�B<����(����Ћ���Q�RLj�j�������QP��(����ҡ���H�A��H���R�Ћ���Q�R��H���P��(���Q�ҡ���P�B<����H����Ћ���Q�RLj�j���8���QP��H����ҡ���H�A��H���R�Ћ���Q�R��H���P��H���Q�ҡ���P�B<����H����Ћ���Q�RLj�j�������QP��H����ҡ���H�A��8���R�Ћ���Q�R��8���P��H���Q�ҡ���P�B<����8����Ћ���Q�RLj�j�������QP��8����ҡ���H�A��X���R�Ћ���Q�R��X���P��8���Q�ҡ���P�B<����X����Ћ���Qj�j���x���Q�RLP��X����ҡ���H�I�U�R��X���P�ы���B�P��X���Q�ҡ���H�A��8���R�Ћ���Q�J��H���P�ы���B�P��H���Q�ҡ���H�A��(���R�Ћ���Q�J��h���P�ы���B�P������Q�ҡ���H�A��8���R�Ћ���Q�J������P�ы���B�P�����Q�ҡ���H�A������R�Ћ���Q�������JP�ы���B�P��x���Q�ҋE����Q��<P�B����W�Ћ���Q�J�E�WP�ыM�����������B�P�����Q�ҡ���H�Aj j������h�cR�Ћ���Q�J������P�ы���B�Pj j�������h�dQ�ҡ���H�A��(���R�Ћ���Q�Jj j���(���h�dP�ы���B�P������Q�҃�@����H�Aj j�������h�dR�ЋF����Q�J$��j0j �|[�j�j ��D8����x����$P�ы���E��B�P������Q�ҡ���H�E��I������RP�ы���B�P��x���Q����F�d8����H�A$��,j0j jj ����h����$R�Ћ���Q�J�E���X���P�ы���B�U��@��X���QR�Ћ���Q�J��h���P�ыF����8�B�P$��,j0j jj ����H����$Q�ҋ�����H�A������R�Ћ���Q�J������PW�ы���B�P��H���Q�ҡ���H�A��X���R�Ћ���Q�R��X���P������Q�ҡ���P�B<��8��X����Ћ���Q�RLj�j�������QP��X����ҡ���H�A������R�Ћ���Q������P��X����RQ�ҡ���P�B<���������Ћ���Q�RLj�j���(���QP�������ҡ���H�A������R�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j���X���QP�������ҡ���H�A������R�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j�������QP�������ҡ���H�A��h���R�Ћ���Q�R��h���P������Q�ҡ���P�B<����h����Ћ���Q�RLj�j�������QP��h����ҡ���H�A�����R�Ћ���Q�R�����P��h���Q�ҡ���P�B<��������Ћ���Q�RLj�j������QP������ҡ���H�I�U�R�����P�ы���B�P�����Q�ҡ���H�A��h���R�Ћ���Q�������JP�ы���B�P������Q�ҡ���H�A������R�Ћ���Q�J��X���P�ы���B�P������Q�ҡ���H�A��X���R�Ћ���Q�J������P�ы���B�P������Q�ҡ���H�A��(���R�Ћ���Q�J������P�ы���B�P�����Q�ҋE����Q��<P�B����W�Ћ���Q�J�E�WP�у��M�������V|�E�<���  ����H�A�U�R�Ћ���Q�Jj j��E�h�cP�ы���B�P�M�Q�ҡ���H�Aj j��U�h�dR�Ћ���Q�J��x���P�ы���B�Pj j���x���h�dQ�ҡ���H�A������R�Ћ���Q�J��@j j�������h�dP�ыF�����j0j �|[	�j���D8�B�P$j ����(����$Q�҉E�����H�A������R�Ћ���Q�M��R������PQ�ҡ���H�A��(���R����F�d8����Q�J$��,j0j jj ��������$P�ы���E��B�P�����Q�ҡ���H�E��I�����RP�ы���B�P�����Q�ҋF�8����H�A$��,j0j jj ���������$R�Ћ���Q�J�������P�ы���B�P�����QW�ҡ���H�A������R�Ћ���Q�J�E�P�ы���B�@�M�Q������R�Ћ���Q�B<��8�M��Ћ���Q�RLj�j������QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j���x���QP�M��ҡ���H�A�U�R�Ћ���Q�E�P�R�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j������QP�M��ҡ���H�A������R�Ћ���Q�R������P�M�Q�ҡ���P�B<���������Ћ���Q�RLj�j��M�QP�������ҡ���H�A�����R�Ћ���Q�R�����P������Q�ҡ���P�B<��������Ћ���Q�RLj�j�������QP������ҡ���H�A��8���R�Ћ���Q�R��8���P�����Q�ҡ���P�B<����8����Ћ���Q�RLj�j��M�QP��8����ҡ���H�I�U�R��8���P�ы���B�P��8���Q�ҡ���H�A�����R�Ћ���Q�J������P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�����Q�ҡ���H�A�����R�Ћ���Q�J������P�ы���B�P������Q�ҡ���H�A��x���R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҋE����Q��<P�B����W�Ћ���Q�J�E�WP�ыM��������E�V|�@�E;E������}�����H�A��x���R�Ћ���Q�Jj j���x���h�dP�ы���B�P�M�Q�ҡ���H�Aj j��U�h�dR�Ћ���v,�Q�J(������VP�ы�����B�P�M�Q�ҡ���H�A�U�RV�Ћ���Q�J������P�ы���B�P�M؃�@Q�ҡ���H�I�U�R�E�P�ы���B�P<���M��ҋ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j���x���QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҡ���H�A��x���R�Ћ]��S�������Q�BV�Ћ���Q�J�E�VP�у��������S����������B�P�M�Q�҃�_^[��]� �������������U���  ����USVWj ��HH��p  h�  R�Ћ���Q�}��j ��h������   j���Ћ���Qj �E����   j���Ћ���Q�J���E�P��d����у�����  �~ ��  ��8����� ������R�ĭ ���ݞ P��8����q ������� ����H�A�U�R�Ћ���Q�Jj j��E�h�dP�у��U�R��8����h
 ����H�A�U�R�Ћ���Q�J�E�P�ы���B�Pj j��M�h�cQ�ҡ���H�A�U�R�Ћ���Q�Jj j��E�h�dP�у�,�U�R�E�P������Q��8���� ��� P�U�R��|���P�YH  ��P�M�Q�LH  ����J�U�RP�A�Ћ���Q�J�E�P�ы���B�P��|���Q�ҡ���H�A�U�R�Ѓ� �������s ����Q�J�E�P�ы���B�P�M�Q�ҋ]����H�Q��S����W�ҡ���H�A�U�WR�Ѓ����Y���S���������8���� ��]����Q�J�E�P�ы���B�Pj j��M�h�cQ�ҡ���H�A�U�R�Ћ���Q�Jj j��E�h�dP�ы�����   �M�Px��(�ҋ�����H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Qj�j�WP�BL�M��Ћ���Q�J�E�P�ы���B�@�M�Q�U�R�Ѓ�����Q�B<�M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҡ���H�Q��S����W�ҡ���H�A�U�WR�Ѓ�������S���1����M�}QWS���Q����}� t��h����ERPWS�����������Q�J��l���P�ы���B�Pj j���l���h�dQ�ҡ���H�A�U�R�Ћ���Q�Jj j��E�h�dP�ы���B�M�@(Q�U�R�Ћ���Q�J�E�E�P�ы���B�U�@�M�QR�Ћ���Q�J�E�P�ы���B�P�M���@Q�ҡ���H�I�U�R�E�P�ы���B�P<���M��ҋ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j���l���QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҡ���H�A��l���R�Ѓ�S���ċ���Q�EP�B�Ћ���Q�E�RP�M�Q�҃����[�������H�A��(���R�E    �Ћ���Q�Jj j���(���hcP�ы���B�P��T���Q�ҡ���H�Aj j���T���hcR�Ѓ�(�} �E    ��  ��d��� �5  �~ �+  ���   �U��� ���   ������   ����Bx�Ћ���Q�R��T���QP�ҡ���P�Rx����(���P��T����҅���  ����H�A�U�R�Ћ���Q�Jj j��E�h�cP�ы���B�P��l���Q�ҡ���H�Aj j���l���h�dR�Ћ���Q�J�E�P�ы���B�@�M�Q��l���R�Ћ���Q�B<��4�M��Ћ���Q�RLj�j���T���QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J��l���P�ы���B�P�M�Q�ҋ���Q��S���ĉEP�B�Ћ���Q�E�RP�M�Q�҃�����������H�I��(���R��T���P�у�����B�P�M�Q�ҡ���H�Aj j��U�h�dR�Ћ���Q�R�E�P�M�Q�ҡ���H�A�U�R�ЋO|�U�� �<� �E    �}  �]�ۍ�    ����H�A�����R�Ћ���Q�Jj j������h�dP�ы���B�P<���M��ҋ���Q�RLj�j������QP�M��ҡ���H�A�����R�ЋG4��N�D����Q�J(P������P�ы���E�B�P�����Q�ҡ���H�E�I�����RP�ы���B�P������Q�ҡ���P�B<���M��Ћ���Qj�j������Q�RLP�M��ҡ���H�A�����R�Ѓ��}� �$  �\ �  ����Q�J�E�P�ы���B�Pj j��M�h�dQ�ҡ���P�B<���M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�ЋGL��N�D����Q�J(P��D���P�ы���E�B�P��|���Q�ҡ���H�E�I��|���RP�ы���B�P��D���Q�ҡ���P�B<���M��Ћ���Qj�j���|���Q�RLP�M��ҡ���H�A��|���R�Ѓ��E�O|�U@���E;�������]����H�A�U�R�Ћ���Q�Jj j��E�h�cP�ы���B�P<���M��ҋ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q��S���ĉEP�B�Ћ���Q�E�RP�M�Q�҃����
����E�O|��U@�E;E��������H�A�U�R�Ћ���Q�Jj j��E�h�dP�ы���B�P��|���Q�ҡ���H�Aj j���|���h�dR�Ћ���Q�E�R(P��D���Q�ҋ�����H�A�U�R�Ћ���Q�J�E�PW�ы���B�P��D���Q�ҡ���H�A�U���@R�Ћ���Q�R�E�P��|���Q�ҡ���P�B<���M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P��|���Q�ҡ���H�A�U�R�Ћ����S�����Q�BW�Ћ���Q�J�E�WP�у��������S����������B�P��T���Q�ҡ���H�A��(���R�Ћ���Q�J�E�P�у�_^[��]� �������������U���   ���SV��H�A�U�WR�Ћ���Q�Jj j��E�h�dP�ы���B�P�M�Q�ҡ���H�I�U�R�EP�ы���B�P<�� �M��ҋ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�ЋM�]��QS��\���R���G�������H�A�U�R�Ћ���Q�Jj j��E�h�cP�ы���B�P�M�Q�ҡ���H�Aj j��U�h�dR�Ћ���Q�J�����P�ы���B�Pj j������h�dQ��݅l�������H�A$��<j0j jj ���������$R�Ћ���Q�J����8���P�ы���B�P��8���QW�ҡ���H�A������R��݅d�������Q�J$��,j0j jj ��������$P�ы����H������BQ�P�ҡ���H�A��H���RW�Ћ���Q�J�����P��݅\�������B�P$��,j0j jj ����d����$Q�ҋ�����H�A��(���R�Ћ���Q�J��(���PW�ы���B�P��d���Q�ҡ���H�A�U�R�Ћ���Q�R�E�P��(���Q�ҡ���P�B<��8�M��Ћ���Q�RLj�j������QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j���H���QP�M��ҡ���H�A��t���R�Ћ���Q�R��t���P�M�Q�ҡ���P�B<����t����Ћ���Q�RLj�j��M�QP��t����ҡ���H�A�U�R�Ћ���Q�R�E�P��t���Q�ҡ���P�B<���M��Ћ���Qj��RLj���8���QP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j��M�QP�M��ҡ���P�B<�M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P��t���Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P��(���Q�ҡ���H�A��H���R�Ћ���Q�J��8���P�ы���B�P�����Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ыU����H��,R�Q����W�ҡ���H�A�U�WR�Ѓ��������Mh�  QS���5������  h�  P������R���)�����������  ������P�M���  P������Q�M��X���R�H� P肪 ����X����d�  �M��\�  ����H�A�U�R�Ћ���Q�Jj j��E�h�dP�ы���B�P�M�Q�ҡ���H�Aj j��U�h eR�Ћ���Q�J�E�P�ы���B�@�M�Q�U�R�Ћ���Q�B<��4�M��Ћ���Qj�j��M�RLQP�M��ҡ���H�A�U�R�Ћ���Q�R�E�P�M�Q�ҡ���P�B<���M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�Jj j�h�c�E�P�у�,��d���R�������}�  ������H�A�U�R�Ћ���Q�J�E�PW�ы���B�P<���M��ҋ���Q�RLj�j��M�QP�M��ҡ���P�B<�M��Ћ���Q�RLj�j��M�QP�M��ҡ���H�A�U�R�Ћ���Q�J��d���P�ы���B�P�M�Q�ҋE����Q��P�B����W�Ћ���Q�J�E�WP�у����������������  ��������  ����B�P�M�Q�ҡ���H�A�UR�Ѓ�_^[��]�$ ����������U����   SV��W�M��z�  ����H�A�U�R�Ћ���Q���   ���E�Pj�M�Q�M�ҋ�����H�A�U�R�Ћ���Q�J�E�PW�ы���B�P�M�Q�҃��E�P��8����n�  ��8���Q�M��o�  ��8������  ����B�P�M�Q�ҡ���H�A�U�R�Ѓ��M�Q�M貆 P�M��I�  �M���  ����B�P�M�Q�ҡ���H�A3�Sj��U�h�dR�Ѓ��M�Q�M��E�  ����B�P�M�Q�҃��E�P�M����  P��� ����Q�J�E�P�у���  h1D4ChCD4C�E���蠢 PSj�U�R����  ��u"�E�P�d�  ���M��]����  3�_^[��]� �]9^�  �N�U����<��H�A�U�R�Ћ���Q�J��t���P�ы���B�Pj j���t���h�cQ�ҡ���H�A��T���R�Ћ���Q�Jj j���T���h\eP�ы�����   �Px��,���ҋء���H�A�U�R�Ћ���Q�R�E�P��T���Q�ҡ���P�B<���M��Ћ���Qj�j�SP�BL�M��Ћ���Q�J�E�P�ы���B�@�M�Q�U�R�Ћ���Q�B<���M��Ћ���Q�RLj�j���t���QP�M��ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J��T���P�ы���B�P��t���Q�ҋE�����Q��P�B����S�Ћ���Q�J�E�SP�у����!�������B�P��d���Q�ҡ���H�Aj j���d���h<eR�Ћ���Q�R�E�P��d���Q�ҡ���H�A��d���R�ЋM�����B�� Q�H����S�ы���B�P�M�SQ�҃���芶��h�  W���}�����tG����H�Q����S�ҡ���H�Qj j�h8eS�ҋE��M��h4  h@  WPQ������h�  W���%�����tI����B�H����S�ы���B�Hj j�h4eS�ыU��E��h�	  hD  WRP���H�������Q�J��D���P�ы���B�Pj j���D���h$eQ�ҡ���H�I�U�R��D���P�ы���B�P��D���Q�ҋE�����Q�� P�B����W�Ћ���Q�J�E�WP�у����@�������B�P�M�Q�ҡ���H�Aj j��U�heR�Ћ���Q�R�E�P�M�Q�ҡ���H�A�U�R�ЋM��� Q����B�H����W�ы���B�P�M�WQ�҃���赴������H�A�U�R�Ћ���Q�Jj j��E�heP�ы���B�@�M�Q�U�R�Ћ���Q�J�E�P�ыU�����H�� R�Q����W�ҡ���H�A�U�WR�Ѓ����+����M�Q�����������B�P�M�Q�ҋE@��;F�E������M���  �E�P�*�  ���M��E�    ��  _^�   [��]� ����������U���  SVW��hG  �������� �K �������������  �������Q�  ����H�A�U�R�Ћ���Q�u���   ���E�Pj�M�Q���ҋ�����H�A�U�R�Ћ���Q�J�E�PW�ы���B�P�M�Q�҃��E�P��\����C�  ��\���Q�������A�  ��\�����  ����B�P�M�Q�ҡ���H�A�U�R�Ѓ���\���Q�M� P��������  ��\����Z�  ����B�P�M�Q�ҡ���H�Aj j��U�h�fR�Ѓ��M�Q��������  ����B�P�M�Q�҃���������  ����H�A�U�R�Ћ���Q���   ���E�Pj�M�Q���ҋ�����H�A�U�R�Ћ���Q�J�E�PW�ы���B�P�M�Q�҃��E�P��\�����  ��\���Q���������  ��\����d�  ����B�P�M�Q�ҡ���H�A�U�R�Ѓ�h�f��\����n�  ��\���Q���������  ��\�����  ��������  ����B�P�M�Q�ҡ���P���   ���E�Pj�M�Q���ҋ�����H�A�U�R�Ћ���Q�J�E�PW�ы���B�P�M�Q�҃��E�P��\�����  ��\���Q�������	�  ��\����n�  ����B�P�M�Q�ҡ���H�A�U�R�Ѓ�h�f��\����x�  ��\���Q���������  ��\�����  �U�R���������  P�֚ ����H�A�U�R�Ѓ��M�Q��������  P譚 ����B�P�M�Q�҃��E�P�������y�  P胚 ����Q�J�E�P����ݕ`�����ݕh�����`�����fRݝp�����x���P������ݕx���Q�荕�����U�Rݝ����������U�ݕ����ݕ����ݕ����ݕ����ݝ�����)  ������   ���   �ҋMj P�E��jx ������   �M����   �Ѕ��  �W�  h1D4ChCD4C�E����s� Pj j������Q���p�  ��uW�U�R�3�  ���3��u����   ���   �U�R�Ѓ��u���������  �������{�  �������p�  3�_^[��]� ����Q�J�E�P�ы���B�Pj j��M�h�cQ�ҋE���P�����M�Q�U�R���������  PW�%  �����H�������H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�ҡ���H�Aj j��U�h�cR�ЋM���Q�����U�R�E�P�������Z�  PW�%  �����ɭ������Q�J�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�Jj j��E�h�cP�ы���B���   �}���j j����W�����M�QP�U�R������PW�$  �����5�������H�A�U�R�Ћ���Q�J�E�P�ы���B���   ��j j���҅�t�E�P����j h�f�ߒ�����ج������Q���   j j���Ѕ�t�M�Q����j hpf訒����衬������B���   j j����P�E�P���N���P�� ����Q�J�E�P�ыM������  ����B�P�M�Q�ҡ���H�Aj j��U�h`fR�Ћ���Q�J�E�P�ы���B�Pj j��M�hXfQ�҃�(�E�P������Q�������i�  P�U�R�E�P�#  ��P�M�Q�#  P�X� ����B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J������P�ы���B�P�M�Q�ҡ���H�A�U�R�Ѓ�$��  h1D4ChCD4C�E��豔 Pj j������Q����  ��u:�U�R�q�  �E�3�P�u��c�  ����u����   ���   �E�P�у��,�������B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�Jj j��E�h4fP�ы���B�@�M�Q�U�R�Ћ���Q�J�E�P�ыU�����H��$R�Q����W�ҡ���H�A�U�WR�Ѓ����d����   3���`���Qǅ`����  ��h�����d�����t�����p�����l����y ����B�P�M�Q�ҡ���H�AWj��U�h�cR�Ћ���Q�J�E�P�ы���B�PWj��M�h$fQ�҃�,�E�P��`���Q������hfR�# P�E�P�M�Q��   ��P�U�R��   ����Q�R�M�QP�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P������Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ыU�����H��(R�Q����W�ҡ���H�A�U�WR�Ѓ������������Q�J�E�P�ы���B�Pj j��M�h�cQ�ҡ���H�A�U�R�Ћ���Q�Jj j��E�h�eP�ы�����(�M�QP������R�O���P�E�P�M�Q�  ��P�U�R�  ����Q�R�M�QP�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P������Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�ыU�����H��(R�Q����W�ҡ���H�A�U�WR�Ѓ���������M�Q���U�������B���   3�Wj���ҋM��{�{������������   ���   ��X����Ѕ���  �ؒ ������   ��X����M����   P�ҋ�������   �B�ω}���=�  �\  ����Q�J��p���P�ы���B�Pj j���p���h�eQ�ҡ�����   �Bx������P��p���Q������R�  P�f� ����H�A������R�Ћ���Q�J��p���P�у��������O�������B�P������Q�ҡ���H�Aj j�������h�eR�Ћ�����   �Bx������P������Q������R�s  P轐 ����H�A������R�Ћ���Q�J������P�у������� ��  ����BH���   ��h�  Q�҃�P��`����l  j��x����_  ��d���3�9�t���~�    @��;�t���|�M��E�    ��� ���}؅���  ������   �B����=�  ��  hF  h�  W��肠�����q  j ���E�   �� ������  h�  W�M�Q���/�������B�P<�M��҅��   V��x�����  �M��R� ������   ���    ������   �B����=)  ��   ������   �Bx���Ћ���Q�Rx�M�Q���҅�us���A� ��T���Q������Rh���3�V�ȉE��� ��tH������F;�T�����������d���I��@;�T���~獅T���P������Q�M�h���V�� ��u�������   �P(���ҋ����(������|���j ��`����0�  ����Q�J�E�P�ы}؃�������   �P(���ҋ��E؅��8�����|����8 ��   ����Q�J�E�P�ы���B�Pj j��M�h�eQ�ҡ�����   ��������R|���E�P�ҡ���H�A�U�R�Ћ����QT3�WP�B�Ѓ�;���  �M�Q����� ����ݕx����U���x����]�Q�B�PHh�  �M��ҋ�|������M���  �}� ��   ������ �E�    ��   3�9s~U��S������ ���   �ȋBx�Ћ�|����U�����������   �Bx�Ћ���Q�ȋBxW�Ѕ�t1F;s|��s��|����U��<���xjjjV���K  ��t�C�<��E�@�E�;������f�������QH�u܋�p  j h�  V�Ћ���QHj ��������p  h�  V�Ћ���QH�����   h�  V��P����Ћ���QH�؋��   h�  V�]��Ћ�X�������(�u�;�t.}+�QV��D����  �jj��+�RQ��D����~  ��X���3���~.�O��]�3�;Q��H�����@�����\���]�;�|ۋ�X���3�3���~��H�����    �@;�|���������\���;�t(}+�PS��������  �jj��+�QP��������  ����BH�P8��P���Q�M��ҋ�   �������������P�����Q������R�?�����݅H����E�    ݅@���݅8���݅0���݅(���݅ ������D  �������u�����   �    �����+�+�+���F�A(��    �������M�݅����������H؋������܅�������H������H���ݝx���݅����H�܅�������H������H����]�݅����H�܅ ������H������H���݅x�����E��\�\������݅����L�H�܅�������H��������ݝx���݅����H�܅�������H���������]�݅����H�܅ ������H��������݅x�����E��Y�Y݅����H܅�������H�����H��������σ�`ݝx���݅����H�܅�������H������H����]�݅����H�܅ ������H������H���݅x����\��E��\��\�������݅����N�H�܅�������H������H����]�݅����H�܅�������H������H����]�݅����H�܅ ������H������H����E�ݝx����E����]�݅x����\��\��E��\�������U�9U���   �M؋������I������D�+�U�+�݅����������H�΃�J܅�������H������H����]�݅����H�܅�������H������H����]�݅����H�܅ ������H������H����E�ݝx����E����]�݅x����\��\��E��\��k�����\����݋��������������;�t&}+�QP�������:  �jj+�PQ�������5  �]�3�3Ʌ��y   ��P�����H������<��� ���u.�r�4��2�� ����t��r��� ����t��r��� ����t���2�4��r��� ����t��r��� ����t���H����A��;�|�����B�M���   j j�҅��a  ����HH�u܋��   j h'  V�ҋ������{  ��\���������;�t,}+�QP�������4  �jj+�PQ�������/  ��\�����(���;�t&}+�QP�������	  �jj+�PQ�������  ����� ��ݕ����3�ݕ����3�ݕ �����P���ݕ���ݕ���ݕ���ݕ ���ݕ(���ݕ0���ݕ8���ݕ@���ݝH������j  ��    ����HD��P����I,������RWP�ы�H����v�Ƀ�Ƀ<��:  ��������8������<����T��@����T��D����T��H����T��L����T��������D�� ������$����P��(����H��,����P��0����H��4����P�������N�I������������P������P������P������P������P�������V�R�Ë�������������X�������X�������X�� ����X������X������4�������F�D�������]������������   ��������� ������$����P��(����P��,����P��0����P��4����P�������D������������P������H������P������H������P�������N�I��������������P�������P�������P�� ����P������P������4�������V�T����������H���4�G;�������M��E�}������SQ�M܍�����RPQW���G���������V����P���   j j���Ѕ�t	������N������萟���ދ������X������   �M����   G��X�����;��3����M��(�  ������ t�{ ~�EVP����������Q�J�E�P�эU�R��  �E�P�E�    ��  ���o  3�Vh�e�������7~��Vh�e�M��)~��������   �M܋Bx�Ѝ�����QP�U�R������P�>  ��P������Q�.  P�x� ����B�P������Q�ҡ���H�A������R�Ћ���Q�J�E�P�ы���B�P������Q�҃� �������J�������H�A�U�R�ЍM�Q��  �U�R�u���  ����u����   ���   �U�R�Ѓ��n������������������Q�J�E�P�эU�R�\�  �E�P�}��P�  ����}����   ���   �E�P�у��}���������B�P�M�Q�ҡ���H�A3�Wj��U�h�eR�Ћ���Q�J�E�P�ы���B�PWj��M�h|eQ�ҡ�����   �Bx��(���Ћ���Q�J���E�P�ы���B�@�M�Q�U�R�Ћ���Q�B<���M��Ћ���Qj�j�VP�BL�M��Ћ���Q�J�E�P�ы���B�@�M�Q�U�R�Ћ���Q�B<���M��Ћ���Q�RLj�j��M�QP�M��ҍE�P�X� ����Q�J�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�у��������3�������B�P�M�Q�ҍE�P��  �M�Q�}���  ����}����   ���   �M�Q�҃��}��U�������Q�J�E�P�ы���B�Pj j��M�hdeQ�ҍE�P� ����Q�J�E�P�у�������R迴 ������   ���   �U�R�Ѓ��������E�    �c�  �������X�  �������M�  _^�   [��]� ���������������VW��3�9>t	V���  ���>�~�~�~�~_^�������������U��Q3�9A~V�u�2@��;A|�^]� ���������������U��EV���
�   ^]� �MW��x/�~;�}(�> t#�~ u%����H��0  h�ch�  �҃�_3�^]� ��;�|���;���_�   ^]� S�;�|�ߋ�+����];���   ^��~�F�I���QP�[��P�c ���N��~�I�ЉV;��'  ������V+ӍR���R��)F+ȍ@��N�N�Q�+�Q�Dc �F����Q���  �@�h�c�h�  �PQ�҃������   �N)^�I[��_�V�   ^]� �V��+Ë^�D�����W�@�Ë]�E;�}-�F+�+�����R��R��R�I��R�b �E��;F}L����Q���  �@�h�c�h�  �PQ�҃����u	[_3�^]� �N�I�ȋE�F�V)^[_�   ^]� ��U��EV���
�   ^]� W�}��x/�N;�}(�> t#�~ u%����H��0  h�ch�  �҃�_3�^]� ��;�|���;���_�   ^]� S�;�|�ً�+����];���   ^��~�F��    QP��R�a ���N��~���V;���   ������V+���R��)F+ȉN�N�Q�+�Q�Va �F����Q���  h�c�h�  �PQ�҃������   �N)^[��_�V�   ^]� �V��+ÍD���~�X�^�A�;�}!�U�F+�+���Q׍�Q��R��` ��;^}C����H���  h�ch�  ��    RP�у����u	[_3�^]� �V���F�^�])^[_�   ^]� ���U�졸��P�B<V���Ћ���Q�M�RLj�j�QP���ҋ�^]� �������������U���VW�}���y
_3�^��]� S�]����  �F��;��ύ�N�U��u(����H��0  h�chA  �҃�[_3�^��]� ��;���  )^�F�b  @����и   +�����ȋF�ڙ�ӉM��ȉE��ډU����������ɋ���]�;�u�;�u�;]�|�;M�r��]�Ù�E�9U��u���;��k����U��N�F�N��F���h�c��u�J�@���  ���hW  R�Ѓ���R�@��hX  �PQ��  �у��ȉ��������F�@�F�щN��~P+Ǎ@���P��+E�Í@��P��@��P�^ �N��ҋ�+E��R�@��RQ�w^ ���  �@���P��+E��@��P�[�a  ��~�V����Q�R�@��R�1^ ���F��@���V�7  �F�D����@����E��F�ʙ�M�;���   	9E���   �E���������ً�����ɋ���]�;������;������;]������	;M�������]�Ù�E�9U������;�������h�c��u'����H�E��@���  ���h|  R�Ѓ��'����Q�M���  �I��h}  �QP�҃��ȉ���Q����F�U��@���N�V�F;�}(�N+Ǎ@���P���P��@��P��\ ���} tG�N;�}"��+��@���R�I�N��j R�[ ���V�[���P���j P�[ ���} tI�N��;�}�F�I�Ћ�+х�t��P�P��Ju�V��ʅ�~��t��P�P��Ku��؋E�F[_�   ^��]� ����U���S�]V���y
^3�[��]� W�}���  �F��;��ˍ9�N�U���u(����H��0  h�chA  �҃�_^3�[��]� ��;��j  )~�F�0  @����и   +�������F�ʙ��߉}����ˋ����ɉE����;�u��E�;�u�;�|�;�r��]�Ù9U�|�;�r��M�F�V��Fы���Vh�c��u����Q���  hW  P�у������RhX  PQ��  �у����� ����V�}�N���F��~@+�ɋ�+U��QӍ��Q��P��Z �F+]��    Q��RP�Z �����P  �ɋ�+U�Q��Q��R�Z ���/  ��~�V��    Q�R��R�hZ ���F����V�  �F�D����@����ȋF����M�;���   ;���   �����ɋ��;��@���;��8���;��0����}�;��#����E�;�����;������h�c��u#����Q���  ��    h|  P�у��"����Jh}  ��    RP��  �Ѓ����������N�]���V�~�F;�} �N�U+���P��P���Q�TY ���} t=�F;�}�N��+���R��j R�-X ���E�V��    Q��j P�X ���M��N_^�   [��]� ����������U�졸��H�QV�uV�ҡ���H�U�AVR�Ћ���Q�B<�����Ћ���Q�M�RLj�j�QP���ҋ�^]���������U��Q�E;�u	�   ]� }+�RP�/���]� jj+�PR�.���]� ����������U��V��W�~��y_3�^]� jjjW�������t�F�M��_�   ^]� ��������f�-\ �����U��M�UV�uW��r�;u��������s��tE��9+�u1��v6�B�y+�u ��v%�B�y+�u��v�B�I+���_��^]�_3�^]�����������U��QV��j �M��I �F���s@�F�M��I ^��]�������U��QVW��j �M��NI �G��t	���sH�G�w����֍M�#��SI _��^��]������f����������U��QW�9��t;j �M���H �G��t	���sH�GV�w����M����I #�t
��j����^_��]�����̰�������������̸   �����������U�������M�P�P�P�P �P(�P0�P8�P@�PH�PP�XX���Q�P�Q�P�Q�P�Q�P�I�H�M��P�Q�P�Q�P �Q�P$�Q�P(�I�H,�M��P0�Q�P4�Q�P8�Q�P<�Q�P@�I�HD�M��PH�Q�PL�Q�PP�Q�PT�Q�PX�I�H\]� �����������U��MV3��� ��t������   ���ȋB(�Ѕ�u��^]� ��������������U���SVW���� �O ���EP�bO P���ʧ �M���  ����Q@�J$�E�PV�ы���B�P4��jh�  �M��ҡ���P�B4jh�  �M��Ћ���E�Q�R8Ph�  �M��ҡ���P�B4jh�  �M��Ћ���Q@�J(j�E�PV�ы]����3��� ��t�d$ ������   ���ȋB(�Ѕ�u�WV���^� ������   �Bj j���ЍM���  ����Q�J�EP�у�_^[��]� �U�졸��U��0SW���HT�Aj R�Ћ؃���u_[��]� V�M�Q��覭 �u���i��   ���   �B�@H�T1 Rh�  �M��Ћ��   ƃ��    ^tH����R��P�B8h�  �M��Ѓ�W�M��ĸ  ����Q�R<�E�Ph�  �M��ҍM��"�  �E�P���G� �M���  _�   [��]� ��U�졸���HSV�ًH�A�U�WR�Ћ���Q�Jj j��E�hcP�ы}���i��   ���   �R�Rx���M�Q��8�   ���������H�A�U�R�Ѓ�����  ����QT�u�Bj	V��3Ƀ��E;�u_^3�[��]� Q�M�M��M�Qh�  �M��[� P��胝 �M���� ������   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   �� P���W� �M�识 ������   �
�E�P�у��u�U�R��身 ����P���   �RH�L8PQh�  �M��ҡ���E�   �E�   �P���   �E�PhT  �M��ҡ�����   ��U�R����   �����    tJ����B�P8�ǐ   Wh�  �M��҃�S�M�袶  ����P�R<�E�Ph�  �M��ҍM���  �E�P���&� �M����  ������   �
�E�P�у�_^�   [��]� ���������U�졸���HSV�ًH�A�U�WR�Ћ���Q�Jj j��E�hcP�ы}���i��   ���   �R�Rx���M�Q��8�   ���������H�A�U�R�Ѓ����H  ����QT�u�BjV��3Ƀ��E;�u_^3�[��]� Q�M�M��M�Qh�  �M��� P���C� �M�軄 ������   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   �ϒ P���� �M��o� ������   �
�E�P�у��u�U�R���z� ��   ���    tK����Q�B8�Ǥ   Wh�  �M��Ѓ�S�M��´  ����Q�R<�E�Ph�  �M��ҍM�� �  �E�P���E� �M���  ������   �
�E�P�у�_^�   [��]� ��������U�졸���HSV�ًH�A�U�WR�Ћ���Q�Jj j��E�hcP�ы}���i��   ���   �R�Rx���M�Q��8�   ���������H�A�U�R�Ѓ�����  ����QT�u�BjV��3Ƀ��E;�u_^3�[��]� Q�M�M��M�Qh�  �M��;� P���c� �M��ۂ ������   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   �� P���7� �M�菂 ������   �
�E�P�у��M�U�R蜧 ���   ل8�   j �5�g�M�Qh  �M��E�   �]�E�]�膐 P���Θ �M��&� ������   ��M�Q����   �����    tK����Q�B8�Ǥ   Wh�  �M��Ѓ�S�M�臲  ����Q�R<�E�Ph�  �M��ҍM���  �M�E�P�	� �M����  ������   �
�E�P�у�_^�   [��]� ������������U�졸���HSV�ًH�A�U�WR�Ћ���Q�Jj j��E�hcP�ы}���i��   ���   �R�Rx���M�Q��8�   ���������H�A�U�R�Ѓ�����  ����QT�u�BjV��3Ƀ��E;�u_^3�[��]� Q�M�M��M�Qh�  �M���� P���#� �M�蛀 ������   �P8�M�Q�҃���uGP�E�Ph�  �M��E�   �E�   诎 P����� �M��O� ������   �
�E�P�у�j �U�Rh�  �M��E�   �E�   �g� P��诖 �M��� ������   ��U�R�Ћu���M�Q���� ���   ǃ��    tJ����Q�   P�B8h�  �M��Ѓ�S�M��Z�  ����Q�R<�E�Ph�  �M��ҍM�踰  �E�P���ݤ �M���  ������   �
�E�P�у�_^�   [��]� U���  ���3ŉE�SVW���SV ��ݕ������\���ݕ������������fPݝ����������Q��0���ݕ����R�荅����ݕ����3�ݝ0���P��P�����h���ݕ����ݕ8���ݕ@���ݕ����ݕ����ݝ������������Q�J��L���P�ы���B�PWj���L���h�hQ�ҍ�L���P�~e ����Q�J��L���P�ы��   ���   +θ����������������d�����  ��p����p����{ �   �}��t{����B�P������Q�ҡ���H�Ij j��U�R������P�ы�\�����������R�C ��`�������H�A������R�Ѓ���`��� t��`���Q�e� ���U�E�RP赼 ������t������j  ����Q���   �J�p�����X���P�ы���B�Pj j���X���VQ�ҡ�����   �R|����X���P���ҡ���H�A��X���R�Ћ���Q�J�� ���P�ы���B�Pj j��� ���h�hQ�ҡ���H�U�I(R��8���P�ы�����B�P��h���Q�ҡ���H�A��h���RV�Ћ���Q�J��8���P�ы���B�P�����Q�ҡ���H�I�����R�� ���P�ы���B�P<��<������ҋ���Q�RLj�j���h���QP������ҍ����P�b ����Q�J�����P�ы���B�P��h���Q�ҡ���H�A�� ���R�Ћ���Q�J�����P�ы���B�Pj j������h�hQ�ҡ���H�U�I(R������P�ы�����B�P������Q�ҡ���H�A������RV�Ћ���Q�J������P�ы���B�P�����Q�ҡ���H�I��@�����R�����P�ы���B�P<��������ҋ���Q�RLj�j�������QP������ҍ����P��` ����Q�J�����P�ы���B�P������Q�ҡ���H�A�����R�Ћ���QH���   j h�  W�Ћ���QHj �E����   h�  W�Ѓ�(�}� ǅx���    ~c3ɋU�t��h���+���|����t+���l����t�+׉��l���+��p�P��|����P��x���B�� ����x���;U�|���t���3�9u���   ��h���݅����݅�����M�݅�����R݅������ҋ��   ��܍h���F����܅P����@܍���������H��� ܍p���܅X����@܍���������H��� ܍x���܅`����@�������H�����Y��Y��Y�;u�|��������؃; �P  �}� �F  ��E�ݕ����Pݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ����ݕ ���ݝ���萘 ��3҃���l���;���  ��x���9U���   ��|����
�d$ ��|����M�t
���   �4v�4�V�t
�4v�4�V�t
�L
�4v�I�4���VR�������Z�����   ������󥋍l������ ����QD��x����R0������QVP�҃�|��� F����x���;u��i�����l�����t���j V���S� ������   �Bj j����j h�  ���ߣ ����   ����Q�J��x���P�ы���B�Pj j���x���h�hQ�ҡ�����   �Bx�����Ћ���Q�J����,���P�ы���B�@��,���Q��x���R�Ћ���Q�B<����,����Ћ���Qj�j�VP�BL��,����Ѝ�,���Q��\ ����B�P��,���Q�ҡ���H�A��x���R�Ѓ��{ ��  ����Q�J��<���P�ы���B�Pj j���<���hcQ�ҋ��   ���   +θ��Q�����������uA����Q��<���P���ĉE�P�B�Ћ���E��Q�JPV�у�W���S����%  �  �����<���R�Q���ĉE�P�B�Ћ���E��Q�JPV�у�W���������   +��   ���Q���������ǅ|���   ����  ǅx����   h)  舔 ����Q�������{  �J������P�ы���B�Pj j�������h�hQ�ҡ���H��|����I(R������P�ы���E��B�P��H���Q�ҡ���H�E��I��H���RP�ы���B�P������Q�ҡ���H�A��L���R�Ћ���Q�R��L���P������Q�ҡ���P�B<��8��L����Ћ���Q�RLj�j���H���QP��L����ҡ���H�I��<���R��L���P�ы���B�P��L���Q�ҡ���H�A��H���R�Ћ���Q�J������P�ы�����   �P|����<���Q���ҋ��E� �E�3���t���9E�~.��I �M���|���9�u�M�P�9� ��t���@��t���;E�|׋�ǅt���    覟 ��t��������   ��t����ȋB(�Ѕ�u㋍t���QV���� ������   �Pj j���ҋ���Q���   �x�����<���P���ĉE�P�B�Ћ���E��Q�JPV�у�W���e������   +��   ��|�����x����   ���Q��������F�|���;��W�������Q�J��<���P�у���\���j j j W���5 ������   �Pj j����3��������������� �������������������Ph�   �������������9Z ������   �M��h����������Jp ���   ���   ��d�����p���x+θ�������������G�d���;��
����   _^[�M�3��< ��]ËJ��<���P�у�3�_^[�M�3��< ��]Í�������o �M�_^3�3�[�e< ��]��������U���SV�񋎤   W���   +ϸ��Q��������3����   �]��E��N �P�-7 ����uAhG  �͌ �����������   ���   M����   �P|Q���ҋN j j W��3 WS������WS���d����~ W��Su�u��������WS������jj��誋 ������   �Bj j���Ћ��   ���   �E��   +ϸ��Q��������C�;��*���_^�   [��]ËB�P�M�Q�ҡ���H�Aj j��U�h iR�ЍM�Q�V ����B�P�M�Q�҃�_^3�[��]�������������U��Q���S�ًH�A�SVR�Ѓ��K$�|�  �K@�t�  �K\�l�  3����   ���   ���   ���   ���   ���   �Cx�C|���   ǃ�   �������   ���   ;�t1�E���;�tW��    �}��E�x����x�   �;�u�_�M����   ���   ���   ;�t/�U�RQPP�V  ���   ���E�P���   QRV��q  �� ���   ^��[��]���������U��QV�񋆈   WP�<�  ���   Q�0�  ���   3���;�t'�U�R���   ���   QRP�yq  ���   P���  �����   ���   ���   ���   ;�t	P�؞  ���N\���   ���   ���   ���  �N@��  �N$��  ����Q�B��V�Ѓ�_^��]�U���D  ���3ŉE�SVW��j�������ˀ  ��,���P�N\�\�  ����Q�Bdj��,����Ћ���Qh�j�x���   h  W�Ћ���Q��jW������P�Bh��,����Ћ�����j@jQ�������@k  ��u%�������J���������������y8 u&���!�������H��������������������j P�ND  �� ��� �  ����Q�J������P�ы���B�Pj j�������h�jQ�ҡ���H�A��t���R�Ћ���Q�Jj j���t���hXfP�у�(��<���R�N\��  ����H�A��d���R�Ћ���Q�R��d���P��t���Q�ҡ���P�B<����d����Ћ���Qj�j�VP�BL��d����Ћ���Q�J��T���P�ы���B�@��T���Q��d���R�Ћ�����Q�B<��T����Ћ���Q�RLj�j�������QP��T����ҍ�T���P�TR ����Q�J��T���P�ы���B�P��d���Q�ҡ���H�A��<���R�Ћ���Q�J��t���P�ы���B�P������Q�ҡ���H�A��,���R�Ѓ���$����
  ��$���Qǅ$���g�b. ��_^3�[�M�3��,6 ��]Ë���B�P��t���Q�ҡ���H�Aj j���t���h�jR�Ћ���Q�J������P�ы���B�Pj j�������h�jQ�҃�(��<���P�N\��  ����Q�J����T���P�ы���B�@��T���Q������R�Ћ���Q�B<����T����Ћ���Qj�j�WP�BL��T����Ћ���Q�J��d���P�ы���B�@��d���Q��T���R�Ћ�����Q�B<��d����Ћ���Q�RLj�j���t���QP��d����ҍ�d���P�OP ����Q�J��d���P�ы���B�P��T���Q�ҡ���H�A��<���R�Ћ���Q�J������P�ы���B�P��t���Q�ҋ������@�����������  �8���ǅ����    �
��$    �I j
��������]  ��Qj h�   ������R�������%e  j������Ph\e��O ������   ������������Q���   ���   �I~  ������R������hxjP�kO ����Q�J������P�ы���B�@j j�������Q������R�Ћ��   ����Q�J�P������P�ы���B�P������Q�ҋ��   ��,Ǆ8�       ��  j������Qhtj��N ����u!���   �D:P������hljQ�N �  j������Rhhj�N ����u!���   �L8Q������h`jR�yN �]  j������PhXj�N ����u!���   �T9R������hLjP�>N �"  j������QhHj�HN ����u-���   ǍH0Q�P(R�� P������h8jP��M ����  j������Qh4j�N ����u-���   ǍHHQ�P@R��8P������h$jP�M ���  j������Qh j�M ����u-���   ǍH`Q�PXR��PP������hjP�lM ���P  j������Qhj�sM ����u-���   ǍHxQ�PpR��hP������h�iP�%M ���	  j������Qh�i�,M ����uZ������R������h�iP��L ��j ������Q��<����
H�����   �����:�   �Q�JP��<���P�э�<����rj������Qh�i�L ����u{������R������h�iP�wL ��j ������Q��t����G�����   �����:�   �Q�JP��t���P�э�t�������B�PQ�ҋ��   Ǆ8�      ���������A�����������������Hr  ��u+�������J���������������y8 u��j P�)<  j��l�����w  �����P�N@�]�  ����Q�Bdj������Ћ���Qh�j�x���   hd  W�Ћ���Q��jW������P�Bh������Ћ�����j@jW��|����Ab  ��u%��l����I��x�����l������y8 u&���!��l����J��������l�����������j P�O;  ������ ����H�A��t���R��  �Ћ���Q�Jj j���t���h�jP�ы���B�P������Q�ҡ���H�Aj j�������hXfR�Ѓ�(��t���Q��T���R�N@��  P������P��d���Q�������P��<���R����P��I ����H�A��<���R�Ћ���Q�J��d���P�ы���B�P��T���Q�ҡ���H�A������R�Ћ���Q�J��t���P�ы���B�P�����Q�҃�(�������v  �������gP�������& ����Q�J��,���P�у���$����wv  ��$���R��$�����% ��_^3�[�M�3��- ��]��Ћ���Q�Jj j���t���h�jP�ы���B�P������Q�ҡ���H�Aj j�������h�jR�Ѓ�(��t���Q��T���R�N@蔔  P������P��d���Q�@�����P��<���R�0���P�zH ����H�A��<���R�Ћ���Q�J��d���P�ы���B�P��T���Q�ҡ���H�A������R�Ћ���Q�J��t���P�ы�l����B��$��x���ǅP���    ��  j
��l����!V  ��Pj h�   ������Q��l����d]  ���   +��   ���Q��������3����   ��L������$    ����Q�J������P�ы���B�@j j�������Q������R�Ћ���B���   �L����@x��������R�Ћ���Q�J���������P�у�Gu2���   +��   ��L����   ���Q��������C�;��X������P���j������Qh�i�)G ������   ��P������   i��   ��:�   P������h�iQ��F ��l����J��j
��l����T  ��Pj h�   ������Q��l���� \  ����B�P��t���Q�ҡ���H�Ij j�������R��t���P�ы��   ����H�A��:�   ��t���WR�Ѝ�t����   j	������Rh�i�HF ������   ��l����Hj
��l����
T  ��Qj h�   ������R��l����M[  ����H�A��d���R�Ћ���Q�Rj j�������P��d���Q�ҋ�P������   i��   ������   �JP�A��d���R�Ѝ�d�������Q�JP�у� ��l����B��x����,�����������|����k  ��u+��l����H��x�����l������y8 u��j P�{5  W�qD �������  ����Q�J��<���P�ы���B�Pj j���<���h�iQ�ҡ���H�A��t���R�Ћ���Q�Jj j���t���hXfP�ы���B�P������Q�ҡ���H�Aj j�������WR�Ћ���Q�J��T���P�ы���B�@��@��T���Q��t���R�Ћ���Q�B<����T����Ћ���Q�RLj�j�������QP��T����ҡ���H�A��d���R�Ћ���Q�R��d���P��T���Q�ҡ���P�B<����d����Ћ���Q�RLj�j���<���QP��d����ҍ�d���P�YC ����Q�J��d���P�ы���B�P��T���Q�ҡ���H�A������R�Ћ���Q�J��t���P�ы���B�P��<���Q�҃�����H�A�����R�Ћ�l����QǄl����i�������� �4i��|���t2������������9u"�������������2�������ȉ
+�������������� t��|�����h  ��|����~5  ��l����B�������g��l����gQ�������� ����B�P��,���Q�ҋ������HǄ�����i���� ��� ������t2�����������9u"������������������ȉ
+������������� t�������Ah  ��������4  �������B��$���������Q��$����2 �M���_^3͸   [��% ��]������������V�������������   ^�����������U���8���3ŉE��M�ES�]VW3�jV�U܈M�R�ˉE؉uȉủu���;  �����uVS�M���s  �u�3��Mȉ�F�F;�t�UȋE̋MЉ�F�N�  �}�;���   �U؋M�R�E�PQW��k  W��   �U�U܋���+�PVS�M��E�   �E�    �E� �/U  �M�Q�M���r  �}�r�U�R�T�  ��j�wV�E�P��� ;  �����u�PV3�S�M��E�   �}��E� ��T  �M�Q�M��r  �}�r�U�R��  ���u؍Eȉ>�~�~;�t�MȋŰEЉ�V�F�"�]�;�t�M؋E�Q�U�RPS��j  S載  ���M�_��^3�[�D$ ��]� ����U���  ���3ŉE�SVW�}��j��������k  j@jW�������V  ��u-�������H������������3ۃ�9Y8u��SP��/  �+�������I��$�����������������j P�/  3�9�P����  ����B�P������Q�ҡ���H�ASj�������h�jR�Ћ���Q�J������P�ы���B�PSj�������hXfQ�ҡ���H�A������R�Ћ���Q�JSj�������WP�ы���B�P������Q�ҡ���H�I��@������R������P�ы���B�P<���������ҋ���Q�RLj�j�������QP�������ҡ���H�A������R�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j�������QP�������ҍ�����P�= ����Q�J������P�ы���B�P������Q�ҡ���H�A������R�Ћ���Q�J������P�ы���B�P������Q�҃���T����nj  ��T���PǅT���g�� ��3�_^[�M�3��! ��]� ����Q�J������P�ы���B�PSj�������h0kQ�ҍ�����P��= ����Q�J������P�ы������B����������  �I j
��������J  ��PSjc������Q�������	R  j������Rh�d�< ����u#���   ���   �F|����+��D�h�D�h�@  j������Ph,k�u< ����u&���   ���   ���   ����+��D�l�D�l�   j������Ph�d�5< ����ue���   ���   @P���   �g  ���   ����+Ћ��   3ɉL�d���   ����+Ћ��   �L�h���   ����+Ћ��   �L�l�  j������Qh(k�; �����c  �Fx�������   �������������������P�@��u�+�P������R�������`S  jj������P��L����
Z  ������r������Q�Մ  ��������������������������R�� �ĉ�x�X�@ �� �܍�L�����C�x3��x�  �;�tPQ��T  ��Q���Dt�;������P�o  ������+�������$I�����������D
���H����   t%��t ~9���   ����+ы��   �L�d�������   ����+Ћ��   �D�d�D�d�������9j  ��L�����F  3ۋ������A�������E����������Z`  ��u)�������H��������������9Y8u��SP�=*  �~|3ɋǺ   ����jSS���P辂  ���;��T  �W�;��K  �H�Q���J�Q��Q�y��4  ����B�P������Q�ҡ���H�AWj�������hkR�Ѝ�����Q�9 ����B�P������Q�ҋ�������;�t*������Q������������RQP��c  ������R蹂  ����L����������������������HǄL���,i��\���ǅ\���,h�K$  ��\����+  ��L����B������ǄL���g�gQ������� ����T����e  ��T���R��T����� ��3�_^[�M�3�� ��]� 3����   �؉��   3ɋǺ   ����jSS���P�1�  ��;�tO;�|��H�Q���O�Q��Q�y����3����   ����H�A������R�Ћ���Q�JSj�������hkP�ы��   R������P��G��P������Q������R����P�g7 ����H�A������R�Ћ���Q�J������P�ы���B�P������Q�ҋ��   +��   ����������������8���  3����   �D8d@3ɺ    ����jj j ���P��  ���   �D9p���   �D8d@3ɺ   ����jj j ���P��  ���   �D9t����B�P������Q�ҡ���H�Aj j�������h�jR�Ћ��   �D8d����Q�J(P������P�ы���������B�P������Q�ҡ���H�������I��@������RP�ы���B�P������Q�ҡ���H�������AR�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j�������QP�������ҍ�����P�5 ����Q�J������P�ы���B�P������Q�ҡ���H�A������R�Ћ��   +��   ��������������Cʃ���x;�� ����������BǄ�����i��P��� ǅ����4it2�������D���9
u"��<�����8����2������ȉ
+���,������L��� t�������B[  ��������'  �������B��T���Ǆ����gQǅT���g�+ �M���_^3͸   [�� ��]� ��U���  ���3ŉE�SV�uW3���j��������������<����������������������������������������V`  j@jV�������6K  ��u$�������H��������������9y8u&���!�������I��������������������WP�F$  9������D  ����B�P��@���Q�ҡ���H�AWj���@���h�jR�Ћ���Q�J������P�ы���B�PWj�������hXfQ�ҡ���H�A��h���R�Ћ���Q�JWj���h���VP�ы���B�P������Q�ҡ���H�I��@������R������P�ы���B�P<���������ҋ���Q�RLj�j���h���QP�������ҡ���H�A������R�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j���@���QP�������ҍ�����P�.2 ����Q�J������P�ы���B�P������Q�ҡ���H�A��h���R�Ћ���Q�J������P�ы���B�P��@���Q�҃���������^  ������Pǅ����g�P ��������;�t*������Q������������RQP�\  ������R�^{  ��3�_^[�M�3��� ��]� ����H�A��P���R�Ћ���Q�Jj j���P���h�jP�ы���B�P��h���Q�ҡ���H�Aj j���h���h�kR�Ћ���Q�J��@���P�ы���B�Pj j���@���VQ�ҡ���H�A������R�Ћ���Q�R��@������P��h���Q�ҡ���P�B<���������Ћ���Q�RLj�j���@���QP�������ҡ���H�A������R�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j���P���QP�������ҍ�����P��/ ����Q�J������P�ы���B�P������Q�ҡ���H�A��@���R�Ћ���Q�J��h���P�ы���B�P��P���Q�ҡ���H�A��d���������3����R��������d�����|����Ћ���Q�J��P���P��x����ы���BVW�P��P���h�kQ�ҍ�P���P�0 ����Q�J��P���P�ы������B��������8���q  ����$    ��d���j
��������<  ��Pj h�   ������Q�������?D  j������Rh�d��. ������   ������P������h�kQ�. ��<�����R��������x  ������P�K\�E}  �������jy  �K\�2|  ������Q�������x  ������R�K\��|  �������6y  �  j������Ph�d�J. ������  ����Q�J��h���P�ы�������������;�t5������RQPP�<X  ��������������P������QRV�X  �� ������������ǅ����   ǅ����    ƅ���� �P���@��u�+�P������P�������E  jj������Q��\����>L  ������r������R�	w  ��������P�� ��3��8�x�   �H�@ �� ��F��\�����H�x�  �;�tPQ�G  ��Q���Dt�>��8���P��a  ����������H�~r�6����Q�J��P���P�ы���B�Pj j���P���VQ�ҡ���H�I��h���R��P���P�ы���B�P��P���Q�ҋ��   +��   ���   ���Q���������� 3��tI3���I ����B��@x��h����R�Ѕ���  �N+���Q��������Gʁ��   ;�r��N+���Q���������LQ���Z  �N+����z���Q���������i��   ��8����OR��h���P�ыN+���Q���������L���x�����\����BǄ\���,i�E�ǅl���,ht��|����R�u  ����|����     �M��    �U��    �E��     �M��    �U��    �E��e���E�    ǅl����g�؅�tN�8��t?j �������c �G��t	���sH�G�w������������g #�t
��j����S�kt  ����p����b	 ��\����H�U�Ǆ\���gR�E�g�� ����H�A��h���R�Ѓ��  ��x��������j������Qh�d�k* ����u7G�������������   +׍�Q������h|kR�������* ���P  j������Ph�d�* ����u5���   �v�ʍHQ�PRP������hlkP��) ��F��d����  j������Qh,k��) ����������ui��|������   �4v���ƍHQPh`kR�u) ���   ƍHQ�PRP������hPkP�S) �苋�   �d1�t1��$��|�����x  jRh(k�H) �����`  ��x������t���   ����+ϋL�t���������������AY  ������P�������J  jj������Q��\����G  ��������5  ������R�� ���     �@   �@    �� �@ ��\�����P�P  ��4���Q�]]  ��H�������X  ������+�������$I�����������t����������[  ���R  �f  ������3�3�3����������������������������������������  �������������   ��$    �������������j/P��@���R�B���P�������[  ��@����W  �������r����P�o( H��������������P�������'G  ��hcW�Y8  ����t*�r�?W�0( ��������HQ��������������F  �������@���������   �D��ы���\$���@�\$� �B�$�Ѓ������������������������������Hk��R����`����$P�҃�`��� ǅ����    �p  ����������+�ɋЋ�����+������ɉ������������� �������r���   �|9p�4��t8�v&�������r���   �������4��|9p�������t������� �������r���   �|9p�4��t�v%�������r���   �������4��|9p�������48������ �������2���   �|9p�4��t�v%�������2���   �������4��|9p�������t������ �������2���   �|9p�4��t�v%�������2���   �������4��|9p�������t������������F�� ��������;�`��������������P�]  ������3���;�t	P��n  ��������������������;�t	S�n  ���������������������  ǅ����   ����  ������ǅ����   �����������������j/P��t���P� ���P��������W  ��t����T  ������+�������$I����������3�������N  �
��$    �I ��������    +�j���j P������ǅ����   ǅ����    ƅ���� �8  ��uP������������s���������������   ����+�P�4��$ �������������ыVp��H�D���   ����   ������������s������j hcP���������u9���������tQ������������s���������������   ����+�P�4��+$ �������������ыVp��H�D�������������r������P��l  ��C;������������������@������;������-�������������   �������xr� ����������������+��������   ��P����# �T3p������+�����H�D:��$I�������������vE��������hcS�O3  ����t*�{r���Ë��������   P�# �T3p��H�D:��������\����HǄ\���,i��l���ǅl���,h�  ��l�����  ��\����B�M�Ǆ\���gQ�E�g�>� ���������������������B�������������������G  ��u+�������H���������������y8 u��j P��  ����Q�J��d���P�ы������BǄ�����i�������� ǅ����4it2������������9
u"�������������2�������ȉ
+�������������� t�������;G  ������ǅ�����g�؅�tN�8��t?j �������2� �G��t	���sH�G�w������������6� #�t
��j����S�:j  ���������1� �������Q������Ǆ����gPǅ����g��� �������� tJ������������;�t+�   ��~r�Q��i  ���^�F    � ��;�uۋ�����R�i  ����������tF������;�t3�   �I �~r�P�i  ���^�F    � ��;�uۋ�����V�_i  ���M�_^3͸   [�� ��]� ����U���  ���3ŉE��ESV��F ����Q���   W�}j j	���Љ����Q���   j j���ЉF����Q���   j j���ЉF����Q���   j j
���ЉF����Q�J������P�ы���B���   ��������Qj������R���Ћ���Q�J�؍�����P�ы���B�P������QS�ҡ���H�A������R�Ћ���Q�FP�������JP�ы���B�P������Q�ҡ���H�A������R�Ћ���Q�J������P�ы���B���   ��$������Qj������R���Ћ���Q�J�؍�����P�ы���B�P������QS�ҡ���H�A������R�Ѓ�������Q�������)h  ������R�N$�*l  �������h  ����H�A������R�Ћ���Q�J������P�у�h�b�������g  ������R�N$��k  �������9h  ����H�A������R�Ћ���Q���   ��������Pj������Q���ҋ�����H�A������R�Ћ���Q�J������PW�ы���B�P������Q�҃�������P�������)g  ������Q�N@�*k  �������g  ����B�P������Q�ҡ���H�A������R�Ѓ�h�k�������f  ������Q�N@��j  �������9g  j�������LH  ������R�N$��g  ����Q�Rhj h�   ������Q���ҡ���H�A������R�Ѓ�j@j������Q��������2  ��u%�������J���������������y8 u&���!�������H�������������������j P��  ��H��� ����Q�J��  ������P�ы���B�Pj j�������h�jQ�ҡ���H�A������R�Ћ���Q�Jj j�������hXfP�у�(������R�N$�f  ����H�A������R�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Qj�j�VP�BL�������Ћ���Q�J������P�ы���B�@������Q������R�Ћ���Q�B<���������Ћ���Q�RLj�j�������QP�������ҍ�����P�� ����Q�J������P�ы���B�P������Q�ҡ���H�A������R�Ћ���Q�J������P�ы���B�P������Q�҃���L�����F  ��L���PǅL���g�� ��_^3�[�M�3���� ��]� ������P�ы���B�Pj j�������h�jQ�ҡ���H�A������R�Ћ���Q�Jj j�������h�kP�у�(������R�N$��d  ������H�A������R�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Qj�j�WP�BL�������Ћ���Q�J������P�ы���B�@������Q������R�Ћ���Q�B<���������Ћ���Q�RLj�j�������QP�������ҍ�����P� ����Q�J������P�ы���B�P������Q�ҡ���H�A������R�Ћ���Q�J������P�ы���B�P������Q�ҋ������H��j
��������%  ��Qj h�   ������R�������-  ��������=  ��u+�������H���������������y8 u��j P��  ������Q�� �������  ����B�P������Q�ҡ���H�Aj j�������h�iR�Ћ���Q�J������P�ы���B�Pj j�������hXfQ�ҡ���H�A������R�Ћ���Q�Rj j�������P������Q�ҡ���H�A������R�Ћ���Q�R��@������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j�������QP�������ҡ���H������R�A�Ћ���Q�R������P������Q�ҡ���P�B<���������Ћ���Q�RLj�j�������QP�������ҍ�����P� ����Q�J������P�ы���B�P������Q�ҡ���H�A������R�Ћ���Q�J������P�ы���B�P������Q�҃�� ������P���~���������Q��������~ t-���   +��   ���Q���������t���T�����������薯��� j h  �e ����L����B  ��L���QǅL���g�_� �M���_^3͸   [�&� ��]� �����̋A �8 t�I0���3���������������̋Q�AH9u�A@V�q<�2�Q ��I0+��^����������������V���F@t�F�Q�^  ���V�    �F �     �N0�    �V�    �F$�     �N4�    �f@��F<    ^������̍Q�Q �Q�Q$�A�A�Q(�Q0�A�A�Q,�Q4�     �A$�     �Q4�    �A�     �Q �    �A0�     ���������U��EVP���� ��f��^]� ���̡��V��H�QV�����V ���   �V(R�V0�V8�V@�VH�VP�VX�V`�Vh�Vp�^x����H�A�Ћ���Q�J���   P�ы���B�P���   Q�ҡ���H�A���   R�Ѓ���^á��V��H�A���   R�Ћ���Q�J���   P�ы���B�P���   Q�ҡ���H�A���   R�Ћ���Q�BV�Ѓ�^��������U�졸�SV��H�QWV�ҡ���H�}�QVW���G�^���   �GS�^�G�F�O �N �W$�V$�G(�F(�O,�N,�W0�V0�G4�F4�O8�N8�W<�V<�G@�F@�OD�ND�WH�VH�GL�FL�OP�NP�WT�VT�GX�FX�O\�N\�W`�V`�Gd�Fd�Oh�Nh�Wl�Vl�Gp�Fp�Ot�Nt�Wx�Vx�G|�F|����Q�B�Ћ���QS���   P�J�ы���B�H���   S�ы���B�P���   SQ��ه�   ٞ�   ����H�Q���   S�ҡ���H�A���   SR�Ћ���Q�B���   S�Ћ���Q�J���   SP�ы��   ��<_���   ��^[]� ��������U��V����f�w� �Et	V�Z  ����^]� ���������U���E��QP�h� ��]� ��������U��S�]V�u;�tW�y�WP�<� �F��;�u�_��^[]� U���E��QP��� ��]� ��������U��S�]V�u;�tW�y�WP��� �F��;�u�_��^[]� U��E]� ������U��E�UV�u��+�QPR�7� ����^]� �������������U��E]� ������U��E�UV�u��+�QPR��� ����^]� ��������������3� �����������U��E���A�I��#���   �} t	j j ��� �   ��t5��� ���EP�M��E�g�� hԱ�M�Q�u��}��E�g�� ��t5�� �UR�M���E�g�E� hԱ�E�P�u��}��E�g�� �� �MQ�M���E�g�� hԱ�U�R�u��}��E�g�P� ��]� ���U��EVP���� ��f��^]� ����U��VW�}W���h� ��g�G�F�O_�N��^]� ������U���SV��W3�WW�~0�~�~�F  �F   �~�~ �~$�~(�~,����jWWj�+W  �؃�;�t9�� ��Q� W�M��E��z� �M��A���s@�A�M��� _�^0^[��]É~0_^[��]����������������U��V���M� �Et	V�iW  ����^]� ���������������U��VW�}W���h� ��g�G�F�O_�N��g��^]� U��V��V�g��� ���Et	V��V  ����^]� �����V����t	P�~� ���    ^�������U���SV��^8�u���g��tMW�;��t<j �M��e� �G��t	���sH�G�w����M����l� #�t
��j���ҋu�S�mV  ��_�N�f� ^[��]�����������̃��d� �������̃��]� �������̃��� ����������3�3������������̃��������������̋�� �����������3���������������� ������������̋A$�8 t�I4���3���������������̋A �8 t�Q0�: ~� � Ë�B�����V���P�҃��u�^ËF0��F ��Q��^����������U���3�S�ىE��E�9E��   	9E��   VW������������|G��tA�E;�|9us�u���C ��UVQR�� u�C0��u�}�)u})0�C 0�(��P���҃��;�t.�MA�E��A��M�U� UU�} �x���|
�} �l���_^�E��U�[��]� ������U���3�S�ىE��E�9E��   	9E��   VW������������|G��tA�E;�|9us�u���E�K$�VPR�� u�C4��u�}�)u})0�C$0�,�E� �P�B���Ѓ��;�t+�   EE��U� MM�} �t���|
�} �h���_^�E��U�[��]� ��U��E��s��s�3ɉP�H�H�H]� ����������U��E��s��s�3ɉP�H�H�H]�  ����������U��A � ��t<�Q;v5�U���t:P�t�A@u"�A0� �A ����t�A ����]� 3�]� ���]� ̋Q V�2��u���^�SW�y0����;�s�_[^��A@u/�A$� ��t&;�w9q<v9A<s�A<�A<�+�I �� _[^�_[���^����������������U��Q�Q$���t9A<s�A<S�]VW����   �A � �E�����   �U��u�Q�A<+�u�]����4��u��u�Q+�u�]������t�5�s��s��]�u���  ����   �A�8�A<+Ǚ;���   |;���   +}��A0�)8�A 8�E��   �A$�8����   �A4� �Q �ǋy$��I4+�   ����   ��E��t|�U��u�Q�A<+�u�]����/��u�Q+�u�]������t�5�s��s��]�u��|8��r2�A�8�A<+Ǚ;�#|;�w+}�A4�)8�I$9��u�]���t�5�s��s�E_3ɉ0^�X�H�H�H[��]� �������U��Q�ES�V��uW�y$���]��t9A<s�A<��s;�u;�s��   �E$tk�A � �E���t_����   ����   �Q�:�A<+Ǚ;�}|;�ww+}��A0�)8�A 8�E$tp�A$�8��tg�A ��A4� ǋy$��I4+�M�E$t?�?�}$��t6��|2��r,�Q�:�A<+Ǚ;�|;�w+}$�A4�)8�I$9���s��s��E_3ɉ0^�X�H�H�H[��]�  ����������U��V�q���Q�F�D�gP� g�[� ���Et	V�O  ����^]� ����U��V�������Et	V�iO  ����^]� ���������������U��V���,h�������h����Et	V�,O  ����^]� ��U��Q�U�E�M���u;AvvSVW�y;�sf+�;�w`�   +���yr�	��E�WQS��� ������t5�U�ERPV�q�������t,�M�+ލ|�WR�^S�� ������u�_^���[��]� �M��yr�	_��^+�[��]� ������U��ASVW�};�s
h(g��� �u+�;�s���]��;�r�Ӄyr�����MRQ�P�ב������u;�s
_^���[]� 3�;���_^[]� ����U��M��3���t>���wjPPQ�2M  ����u(�EP�M��E    �D� h���M�Q�E��f�� ��]� ������������̋A �8 t�Q0�: ~����I ��P�� Ë�P���������U��}�Q�Q�Q�Q �Q�Q$���AP�Q(�Q0�AI �A�A�Q,�Q4�     �A$�     �Q4�    �A�     �Q �    �A0�     �E��t�P�Q�Q�P�A �A$�Q0�Q4�AT����QL�AD    ]� ��U��E��u�yr�	�E�U�]� �yr�	MP�EPQ�I� ��]� ��U��QV��W�N��g�e� jj j j�K  ������t0S�*� ���� j �M����� �C���s@�C�M��� [�3��~8�F�F�N�N �V�V$�F�F�N(�N0�V,�V4�     �F$�     �N4�    �V�    �F �     �N0_���    ^��]�U��ES�]V���F<    �F@����   ��<tyWS�ND�������ESPW�� ���F@��F<u�N�9�V �:�N0��N@��u7��u�ǋV�:�N$���+ЋF4Ӊ�N �9 u�V�:�F �     �N0�9�N@_^[]� �����������U��M��3���tN��"""wjPP����+����P�BJ  ����u(�MQ�M��E    �T� h���U�R�E��f�� ��]� �������������U��M��3���tG���Gwi��   jPPQ��I  ����u(�EP�M��E    ��� h���M�Q�E��f�1� ��]� ����U��M��3���tN��I�$	wjPP��    +���P�rI  ����u(�MQ�M��E    �� h���U�R�E��f��� ��]� �������������U��M��3���tH�����?wjPP��    P�I  ����u(�MQ�M��E    �� h���U�R�E��f�`� ��]� ���U��E�M�U ��E��   ]� ����U��E�M��   ]� ������������U��E+E�M;�s��]� ����������U���EV����ft	V�I  ����^]� ��������������U��ES�];��c  VW�}�p��    ����H�A�V�WR���F��_��_�N�O�V�W �F�G$�N�O(�V�W,�F�G0�N �O4�V$�W8�F(�G<�N,�O@�V0�WD�F4�GH�N8�OL�V<�WP�F@�GT�ND�OX�VH�W\�FL�G`�NP�Od�VT�Wh�FX�Gl�N\�Op�V`�Wt�Fd�Gx�Nh�O|����B�@���   Q�VlR�Ћ���Q�R���   P�N|Q��ن�   ٟ�   ����H�I���   R���   P�ы���B�@���   Q���   R�Ћ��   ���   ���   �V��(���   ;��������_^[]ËE[]������U���SV3�S���� �E�^�^�^�^�^�^�^�^ ;�u(�EP�M��E�h�� hL��M�Q�E��f��� PV��� ����^[��]� ���V��WV�_� �F3���;�t	P�� ���~�F;�t	P�n� ���~�F;�t	P�[� ���~�F;�t	P�H� ���~_��^�� ������������U���8SW�}3ۉ]���tz9uvVjSSj�E  ������tO�E� �H�   ��u�HQ�M�������M�Q�F    �Xg�6� ��V�H�N�P�V�@���F�3��7^��t�M�����_�   [��]��������U��V��F�Xg��~�FP�q� �y�NQ��E  ���E��ft	V�E  ����^]� ��������U��U��t�Ay8 u���URP�.���]� ����������V��F � ��t;�N0�	��~�F0��v �@�� ^Å�t�V0�: ~����F ��Q���	��P���҃��u�^ËF �8 t�N0�9 ~��^Ë�P��^��������U���V���F@Wt �~$���t�N<;�s�F4� +��N4��E���u
_3�^��]� �V$�:S��t�N4����;�s�	�-  �F@u=��u3���F4�N�+ߋ���� s�    ���t������+�;�s��u��u[_���^��]� �P�ND�E��3������F��U���tSRW�� �U�����u0�N�~<�9�F$�8�N4�E���F@uE�F�8�N �9�F0�    �e�F$��+�N<� �N��+�+��N$ǉ��+�M��F4��F@t�N�9�F �     �N0�9� �F$��F � �^+�ǉ;�~ +ȉ�F0A��F@t	R�rC  ���F4�N@��E�v$�[�Q�_�^��]� ��������������U��V��F�MW;�s
h(g�� �}+�;�s����tP�VS��r���ރ�r����+��P��SR�� �F��+ǃ~�F[r�� _��^]� ��� _��^]� ��������������U��E�MPQ�� 3҃������]��̋AT��tP�� Y�̋AT��tP�� Y��V��~T t#��Pj��҃��t�FTP��� ����y���^�3�^ËQV�2�AH;�t�q<�q0�6W�y 7_�q@��Q ���+ЋA0��I�^�������������U��S�]V��F � ��t-�N9s&���t�P�;�u�F0� �v ��C���^#�[]� �FT��t8���t3�~D uP��P�� �����u�N �FH9t�Έ�I���^��[]� ^���[]� ��������V��F ���t�V0����;�s�^Ë�PW���ҋ����u_�^Ë�PW���ҋ�_^��������������U��W���OT��t@�UV�u��u��Eu�   �3�VPRQ��� ��^��u�OTjQ���j�����_]� 3�_]� ������������U��j�h`Pd�    P��SVW���3�P�E�d�    �e���u�E�������v���'�^���鸫�������;�v�����+�;؍<v������E�    �OQ�N�E����؉]��E������3�e��E�E�E�@P�M�������E��E�   ��Ëu�}�]�M��t�~r����QPS�i� ���M�~r�R��?  ���M� ��~�N��r��� �M�d�    Y_^[��]� �u�~r�P�?  ���F   �F    � j j �N� �������U���j �M�� � �=l� ����E�u+j �M��� �=l� u�h�@�h��l��M��� S�]�VW�=l�;xs\�H�4�����   �x t�� ;xs
�P�4���uh�u���ua�E�SP�H��������uhpi�M��� h���M�Q�� 3�뮋u�j �M�5���^� �F���s@�F�M�r� V�� ���M��a� _��^[��]�U��M�E+�V���4�    �EVQP��� ���^]� �����U���(SW�}3ۉ]���tW9uSVjSSj�l=  ������t,�E� �H�   ��u�HQ�M������F    �lh�3��7^��t�M������_�   [��]�����������U��W�}��tV�u�   �^_]�������U��M��t	�EP�=���]������������U��j�h�Pd�    PQSVW���3�P�E�d�    �e��E�    �]�}�u��$    ;utVWS�s�������x�}��x�u���E������ǋM�d�    Y_^[��]�j j ��� �������������̋V�qX�H�D1�,iW�N��F�,h�����N�������V��B�D0�gV�g�k� ��_^��������V��~r�P�<  ���F   �F    � ^����������V���@W3��D0u�D08��ȋB4�Ѓ��u�   ��I΅�t�Aǃy8 u��j P�����_��^��U��S�Y���HV�sX�D1�,iW�N��F�,h������N�� ����V��B�D0�gV�g�� ���Et	S��;  ��_^��[]� �����������U����A0SVW�8j �M��}��U� �G���s@�G�M��i� �M�Q������j �M����)� �G��t	���sH�G�w����M����0� #�t
��j���Ћ�E�RP����_^[��]� ����U��j�h�Pd�    P��SVW���3�P�E�d�    �e���u��H΋A���  �I<��t�b����} ��   ��B�L0��t�D00�8�}j �M��g� �G���s@�G�M��{� �MQ���������M�-���E�    ��B�L08�����E���uj j��I�������ЋG�PHu*�E�������I΃y ue��M�d�    Y_^[��]� ��Q�L28����렋M��@��H���x8 u�����H�Hu�E�������$Ëu��j j �� �A���y8 u��j P�b���2��M�d�    Y_^[��]� ������������U��j�h�Pd�    P��SVW���3�P�E�d�    �e���E=���?v
h@g�m� �N+��;�sSP�N�Z����؉]��E�    S�VR�P�������E�������~+�����t	P�9  ���M���V���F��M�d�    Y_^[��]� �M�Q��8  ��j j �� �������U��U��V�p�d$ �@��u��M+�P�ARPj �'��������^]���������������U���j �M��0� �=�� ����E�u+j �M��� �=�� u�h�@�h�����M��� S�]�VW�=��;xs\�H�4�����   �x t�� ;xs
�P�4���uh�u���ua�E�SP���������uhpi�M��� h���M�Q�� 3�뮋u�j �M�5���n� �F���s@�F�M�� V�� ���M��q� _��^[��]�U��j�h�Pd�    P��|SVW���3�P�E�d�    �e��E�    �]�}�u��I ��t-jxj ��x���P��� ��x���QVS�^�����O�}��x�u���E������M�d�    Y_^[��]�j j ��� �������������U��j�h Qd�    P��SVW���3�P�E�d�    �e��}�}��E�    �]�u��;utVWS����������   �}���   �u���E������ǋM�d�    Y_^[��]Ëu�};�t��$    ���������   ;�u�j j �� ������U��EVWP����������B�����Є�t�GD    _^]� �ωwD�'���_^]� �U��S�]V��F���+�;�w
hg��� ��t|W�<���v
hg��� �N;�s5PW���������tT�U�FRSP��������~�~r5��8 _��^[]� ��uԉ~��r�_�  ��^[]� _��^�  []� ���8 _��^[]� ��������U��S�]V��MW�y;�s
h(g�� �E+�;�s��;�uj��W�������Sj ������_��^[]� ���v
hg�� �F;�s(�FPW�������M��th�   9Ar�	9Fr*��(��u�~��r�_�  ��^[]� _��^�  []� ��W�QP�� ���~�~r��8 _��^[]� ���8 _��^[]� ���������U��j�h Qd�    P��SVW���3�P�E�d�    �e���u�3ۉ]�^�^�u܋�H�L18;�t��B��j���������tw�}��|p�]��td�E�    ��Q�L28�����E���u�M��:�M;�u�F�V ��H�L18� ��������]����}��u|��uo�M��E������]�E�  �NNu���Ӌ�H΅�t�Ay8 u��j P������E܋�Q�L8��t��P�ҋƋM�d�    Y_^[��]� �F�V �M�A�M��B�L08�����)����M��B��H���x8 u�����H�Hu�E�������+Ëu��?���j j �� ���U��V��~T ��   �E�M�UPQR�� ����t}WjP�������F8�8j �M�}�+� �G���s@�G�M�?� �MQ���������B�����Є�t�M�FD    ��v��_��^]� �Ή~D�K����M��v��_��^]� 3�^]� ����U��A�UV�1W+ƿ���?��+�;�s
h@g��� Q+���;�v!�������?+�;�s3���;�s��R����_^]� ����U��S�]V���tY�N��r����;�rG��r���ƋV�;�v3��r��MQ+�SV������^[]� �M��Q+�SV�������^[]� W�}���v
hg�D� �F;�s�VRW���S�����t[�~r*��(��u�~��r�_�  ��^[]� _��^�  []� ��WSP�U� ���~�~r��8 _��^[]� ���8 _��^[]� �����������U��E�UP�Ej ��Q�MQRP������]� �����������U��j�h@Qd�    P���   SVW���3�P�E�d�    �e��}�}��E�    �]�u��t0��$��������PWS�x�������$����J���N�u���   �}���E������M�d�    Y_^[��]Ëu�};�t���������   ;�u�j j �� ��������������U��j�h`Qd�    P��4SVW���3�P�E�d�    �e�3��}��E� �u�u���H�L18��t��B��j ���9�������   ��A�D00��]�j �M���� �C���s@�C�M��� �U�R�������E�j �M��̼ �C��t	���sH�C�{����׍M��Ӽ #�t
�j�ϋ��j�j �]�������E�    ��P�D2 �L2$��|��t�EЉMԃ��s�EȉM����������}؋L28������E���t	���uo�M��E������}��@3ۉ\0 �\0$8]�u����I�;�t�A�9Y8u��SP������E���J�L8;�t��B�ЋƋM�d�    Y_^[��]��ЋM܋I�QHu�Pj�������E�O�}؋�B�L08�q����Q����M��B��H���x8 u�����H�Hu�E������1Ëu�/���j j �q� ����������U��EW�};�tsV���   ����H�A�VR�Ћ���Q�BV�Ћ���Q�J�F�P�ы���B�P�N�Q�ҡ���H�A��\���R�Ё��   ��\�����;�u�^_]�������������U���,���3ŉE�V��F 3�9t.�N0� �	�;�s!�F0��v ��P�� ^�M�3��T� ��]�9VTu���^�M�3��=� ��]ËN�FHW9u�F@�~<�9�N ��N0+��9VDu7�vTV�� �����t_��^�M�3���� ��]�_���^�M�3���� ��]ÉU��U��VTSR�E�   �P� �������   �Pj�M��%����M�E��Ѓ�s�U���U��ND�9�]�S�]�S�]�S�]�SRP�FLP�G�Ѕ���   ��~G��u{�}�r`�}��E�s�E�jP�M�jQ�� �u߃��M������[_��^�M�3��*� ��]ÍM�9M�uM�}��E�s�E��U�+�Rj �M��(����FTP�� ������3����M�����[_���^�M�3���� ��]Ã}��}�s�}�+}�}���~��E؋VT�L�ORQ�� ������uߍM��Z����M�[_��3�^�� ��]��������U��QS3�VW���]�9]t�|i�GXg��H�g��_�_�r��������Gj �ΉF8�^<������F@9^8u�F��SP���'�����H�]�,i�O�������3��G,h��u�   ��u����t����t���M�y�Qr�	PRQ�O�I�����_^[��]� ��������������U��V��FW�};�s1�;�w++���;Fu	j��������F��t*�����F_^]� ;Fu	j�������F��t���F_^]� �����������U���$���3ŉE�SW��3�9_D�  8_I�  ��Pj��҃��u_2�[�M�3���� ��]ù   3��]��M�E��E��E�   ��s�E��XV�E��]�Ѓ�s�U���U��OD�1�]�SRP�GLP�F�Ѓ� t#Ht$���M�t{�D���^_2�[�M�3��o� ��]��GI �]�E��ȃ�s�M��u�+�t"��s�E��OTQVjP�A� ��;�u$�]�E��I t���j���Vj�M������T����M�눍M������^_�[�M�3���� ��]ËM�_3Ͱ[��� ��]�����U��E�UP�Ej ��Q�MQRP�B�����]� �����������U��UV���W�F   �F    � �x�@��u�+�PR���>���_��^]� ������U���,���3ŉE�S�]3�V������  �V$W9t0�N4��9�;�s#�	�v$��H_��^��[�M�3��� ��]� 9FT��  �V�NH9
u�N@�~<�:�V �
�V0+ɉ
9FDu.�vT��VP�T� ������i  _^��[�M�3��� ��]� �   �ЈE��]܉M�U��E��E�   ��s�U��B�E��]�Ѓ�s�U���U��ND�9�]�SRP�U�R�E�P�U�R�FLP�G�Ѕ���   ��k�]�E��ȃ�s�M��}�+�t&��s�E��NTQWjP�&� ��;���   �]�E��U��FI9U�u{���s����}� �M���   Wj�\����S�����ur�FT�M�PQ��������t �u�M�����_��^[�M�3��� ��]� �M�����c���_��^[�M�3��� ��]� �M��F����E_^[�M�3��p� ��]� �M��(������_�M�^3�[�R� ��]� ��U��SV��N �FHW9u�}u�~D u�]�}��������}�]�~T ��   ���������t}���u�}t�E�NTPWSQ�_� ����u[�FT�URP�T� ����uG�N�FH9u�V<�F@��N ��V0+���E�M�U_�H�NL^�     �@    �P�H[]� �E��s��s_�H3�^��H�H�H[]� ������U����ES�]V��M�M�3�W�}�E�9NT��   ��������tz�FT�U�RP�� ����uf���t�VTjSWR�w� ����uL�NT�E�PQ�l� ����u8�U�ΉVL������E�M��U�_�H�NL^�     �@    �P�H[��]�  3ɋE��s_���s^�P�H�H�H[��]�  �����������U��VW�}��;�t`�~r�P��#  ���F   �F    � �s�OAQWV�N� ���
���    �G�F�O�N�G   �G    � _��^]� ����������SV��3�W��9^Tt������u3��FTP�v� ����t3��N�N�^P�^I�V�V �N�N$�F�F�V(�V0�N,�N4��V$��F4��N��V ��F0��^T�����_�^D�NL^[������������U��j�h�Qd�    P��SVW���3�P�E�d�    �e���}��"""v
h@g謵 �N+���������������;�srW�N�I����E��E�    P�NQ�R�������E�������N+˸����������������t	S�%"  ���E����+ȋE�ȉV����+ύȉV��M�d�    Y_^[��]� �E�P��!  ��j j �� �������U��V�u�~r�P�!  ���F   �F    � ^]�����U��EV���F�@   �@    �  ���t#PQ�������Q���D��t�    ^]� ��^]� �U��V��~T �4it�N�FH9u�V<�F@��N ��V0+���~P t���������<����Et	V� !  ����^]� ������U��S�V�q+󸉈����E��������"""+�W;�s
h@g�ֳ �y�+����������������;�v!����"""+�;�s3���;�s��P����_^[]� ��U��j�h�Qd�    P��SVW���3�P�E�d�    �e���}���Gv
h@g�L� �N+���Q���������;���   �NW�W����E��E�    P�NQ�R�������E������N�+˸��Q�����������t�EP�FP�FPS�)����Q�  ���Ei��   �M���Fi��   ��~��M�d�    Y_^[��]� �U�R�s  ��j j �>� �������U��V�u;utoSW�}3�;�tR�r�P�;  ���G   �_��~s�NAQVW�ʺ �������F�G�N�O�F   �^�����;uu���_[^]ËE^]����������������U��V�uW�};�t*��~r�P�  ���F   �F    � ��;�u�_^]����U��QSV�u��W�{��+��������������}�;�vE�����+΍�;���   ��;���   ��I ������x�   ��x�;E�u�_^�S[��]� si��+�R��� ����E�{Pj �KQ��+���������������j +�QW�_����{��+���������������+�������+΍ωS_^[��]� ����������U��QS3�VW�ىE�9Et��i�Chg��Q�g�C�C��x����@����sj �ωw8�G<    �����8 �G@u�G��j P���������Q����i�����N�N �4i�FP �FI �F�F�V�V$�N(�N03ɍF�F�V,�V4��F$��V4�
�F��V �
�F0��NT���_�VL�ND^��[��]� ����̋A��PV�q��D
��i�~T �4it�N�FH9u�V<�F@��N ��V0+���~P t�������������F��H�D1�g^�U��QVW�9+׸��Q��E��������G+�;�s
h@g�9� �Q�+׸��Q���������;�v!�����G+�;�s3���;�s��P�n���_^]� ��������U��M��t�E�A   �A    P� �����]�����������U��j�h�Qd�    P��SVW���3�P�E�d�    �e��}�}��E�    �]�u��;utVWS���������}���u���E������ǋM�d�    Y_^[��]Ëu�};�t�]VS�C�������;�u�j j �׿ ����������������U��SV�uW���_��+���Q���������;�v=i��   7;���   �EPVSS�����MQ���G�WRPV�	����� �w_^[]� sc��+�Q���.����U�_Rj �GP��+���Q��������ʋ�j +�RS������_��+���Q���������+�i��   ���w_^[]� U��VW�y��wh���^���V�g��� ���Et	W��  ����_^]� ��������U��E�UP�Ej ��Q�MQRP�"�����]� �����������U��QV����t�M�Q�N�VRQP������R�  ���    �F    �F    ^��]��������������U��QV��F�;�t(�U�WRQPP������V���E�P�NQRW�_����� �~_^��]����U��j�h�Qd�    P��SVW���3�P�E�d�    �e���}��I�$	v
h@g��� �N+��$I�����������;���   �NW�e����E��E�    P�NQ�R�������E������N�+˸�$I�������������t�EP�FP�FPS�����Q�]  ���E��    +ЋE���N��    +׍��N��M�d�    Y_^[��]� �U�R�  ��j j �� �����������U��S�V�q+�$I���E��������I�$	+�W;�s
h@g�� �y�+���$I�����������;�v!����I�$	+�;�s3���;�s��P�i���_^[]� ��U��V�uW���O;�sA�;�w;+�$I�����������;Ou	j���F������    +ƍ��O��t/P�;Ou	j��� ����O��tV�A   �A    � �"����G_^]� ��������U��V�uW���O;�sE�;�w?+�$I�����������;Ou	j���������    +ƍ��O��t7j�j P�;Ou	j�������O��tj�j V�A   �A    � �*����G_^]� U��VW�}��;�tG�S3�;�t�MQ�N�VRQP�g����R�/  ����^�^���O�N�W�V��_�_[_��^]� ���U��EW�};E,t<��MQ�ML������E��t#�URP�#�����Q���Dt3��E��E;E,uŃ}$�EL�r�MQ�  ���}D�E$   �E     �E r�U0R�}  ����_]������U��Q�ML�E��U,SV�uPQ�� �ĉ�H3�j�S�E0�A   �YP�������M�� �ĉj��HS�U�A   �YR������V������L�}$r�EP��  ���}D�E$   �] �]r�M0Q��  ����^[��]��U���(�ML�E�U,SVWQ3�j��E�S�E0�   P�M��U܉u�]��]��X����M܃� �ĉj��HS�U��q�YR��7����   9}�r�E�P�d  ���Mj�S�U�M�R�M��u�]��]������M܃� �ĉj��HS�U��q�YR������9}�r�E�P�  ���M�Q����� �U���H�EL�9}$r�EP��  ���u$�] �]9}Dr�M0Q��  ���E�_^[��]�������U�조���t]��]���������������̡�����   ���ǀ�   �J�p   �������������������������������U��E�� tHt3�]ù���O �����]ø   ]������j j j jdjdhZ� j���>  � ����U���VWjhHljjH�H  ������t���(T �N�l�
����3�����H�A�U�R�Ћ���Q�Jj j��E�h8lP�у��U�R�M��kZ �8Vj�AD ��PWj j�3D ��PhZ� �eV ���M����X[ ����H�A�U�R�Ѓ�_��^��]�������������U��V��N�������{S �Et	V�  ����^]� �����U���EV����lt	V�h�������^]� ��������������U��U�BV�uW�}�g��'���F�g��'��������������AzT�M�B�f��&���A�f��&����������u.��!�B�a����!�G�a����������u_�   ^]� ��_3�^]� �������������U��M��t	��Pj��]������������U����QT��+QP����*��S��VW�����3҉M��w���|{�IP�4v���(   �+ٍA �]���]���H��D�r�H��u�4����_���`���@��H��@��H������@��H��@��H������@��H��@��H�����;�|��M��u�;�}1�YP�R��v�����+��D���L�ȃ�O����u���l_^[��]�����U����US�]VW���M���GP���R�4ЋU���R�Ѝ[�D����f�E���U��&���B�f� �&�����_����z_^2�[��]� 3�9]~9;]t.;]t);]t$���OP�@���M�PQRV��������u��M�U�C;]|�_^�[��]� ����������U���S�ًKT+KP����*����V�����]���D  3ɋƺ   ����W���Q�z��������ˉ}��E� �������c����Au3���~$�d$ ��@;�|��3���~�N���@I;�|��E��ƉE��6�^�����  �u���$    �E��M�]��I�M����  ;�3ۍK�M;��E    �}G9}�3��E��M��UPQ�M�WRS�A������Q  �}� �E��M�����<��F�U�M��  �]�;�s.��U�;�w%��+���;Fu	j���B  �F��t �����;Fu	j���$  �F��t��F�F�M�U�M�;�s+�;�w%��+���;Fu	j����  �F��t#�����;Fu	j����  �F��t�M��F�F�U�}�;�s2�;�w,��+���;Fu	j���  �F���$  �����  ;Fu	j���q  �F����   �8��   �}�;�s.��U�;�w%��+���;Fu	j���:  �F��t �����;Fu	j���  �F��t�8�F�F�M�U�M�;�s+�;�w%��+���;Fu	j����  �F��t#�����;Fu	j����  �F��t�M��F�F�U�]�;�s+�;�w%��+���;Fu	j���  �F��t �����;Fu	j���p  �F��t��E�M��F@;�}�U���I �<��|��@;�|�I�	�M��E���M����L����}�W�s�����_^[��]� �������U��]�w���������̋�3�� �l�H@�HD�HH�HP�HT�HX�H`�Hd�Hh�����������V��W��l�F`3�;�t	P�������~`�~d�~h�FP;�t	P�������~P�~T�~X�F@;�t	P�ռ�����~@�~D�~H_��l^�jp虼��3Ƀ�;�t"� �l�H@�HD�HH�HP�HT�HX�H`�Hd�Hh�3�������������U��M��3���tD�����?w��    P�<�������u(�MQ�M��E    �N� h���U�R�E��f蔯 ��]� �������U��j�h Rd�    P��SVW���3�P�E�d�    �e���E=���?v
h@g荝 �N+��;�sSP�N�J����؉]��E�    S�VR�P��������E�������~+�����t	P蔻�����M���V���F��M�d�    Y_^[��]� �M�Q�c�����j j 辮 �������U��A�UV�1W+ƿ���?��+�;�s
h@g�ל Q+���;�v!�������?+�;�s3���;�s��R�����_^]� ����U���E��P���\$�E�\$�E�$��]� �����������U��E�I@�U�@�����M��@�U��@�]� �����U��E�I@�U�@�����M��@�U��@�]� �����U��M��3���tF�����
w�I���P��������u(�MQ�M��E    �,� h���U�R�E��f�r� ��]� �����U��M�U�E;�t.V�1�0�q�p�q�p�q�p�q�p�q�p����;�u�^]�U��E��t%�M���Q�P�Q�P�Q�P�Q�P�I�H]����������������U��j�h Rd�    PQSVW���3�P�E�d�    �e��E�    �]�}�u��$    ;utVWS�s��������}���u���E������ǋM�d�    Y_^[��]�j j �e� ��������������U��E�UP�Ej ��Q�MQRP�R�����]� �����������U��j�h@Rd�    P��SVW���3�P�E�d�    �e���}�����
v
h@g�,� �N+����*���������;�shW�N������E��E�    P�NQ�R���R����E�������N+˸���*�����������t	S�������E�@�E�ȉV��ȉV��M�d�    Y_^[��]� �E�P�߷����j j �:� ���U��QVW�9+׸���*��E������򺪪�
+�;�s
h@g�I� �Q�+׸���*���������;�v!���꿪��
+�;�s3���;�s��P����_^]� ��������U��QV��FD�N@W;�t�U�RQPP�2������FD�FT�NP;�t�U�RQPP�������FT�Nd�~`;�t ��+�S����    SQW�/� ��߉^d[_^��]�U��V�uW���O;�sb�;�w\+𸫪�*���������;Ou	j���������v���G��tc���Q�P�Q�P�Q�P�Q�P�I�H�G_^]� ;Ou	j�������G��t"���N�H�V�P�N�H�V�P�N�H�G_^]� ������������U����E�A@���Q@�U��E���U��E���U�;Bu+���������Q�Y(�Q�Y0�Q �Y8�M�Q���������]� �������A������Au���Q���Q����z�Q�A ������Au���Q ���A(������z���Y(����A0������z���Y0����Q8����A�{����M���Q���n�����]� ��������U����EV��M3���^�V@�u�;VD�n  �FT�NP;�t�URQPP�������FT�F(S�fW�F0�f�F8�f ��������Au%������Au��3�������Au�Y�]�   �_��X������z+��������Au$�ع   ������Au3��Y�-�   3��$��������ٹ   ����z3��Y��3ۿ   �VD+V@����*���������ЋF@t;�؍<��4ȉU��M��]�E��P�]��P��]��;����������Muԋu��Nd�^`�~`;�t!��+�����PQS�E�'� �M��ˉOW��������W+���������E��t�_[^��]� _3�[^��]� ������U��V���u����Et	V艳������^]� ��%`�%`�%`�%`������U��V�u���t����QP��Ѓ��    ^]���������̡���H��@  hﾭ���Y����������U��E��t����QP��@  �Ѓ�]����������������U�졸��H���  ]��������������U�졸��H��  ]�������������̡���H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�Ѻ ������u_^]Ã} tWj V�|� �������_�F���   ^]���U�����E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]Ã�s�   VW�xW�(� ������u_^]À} tWj V�Ӛ �������_�F���   ^]����������U��M��t-�=�� t�y���A�uP�{� ��]á���P�Q�Ѓ�]��������U��E���� ]�̡��V��H�QV�ҡ���H$�QDV�҃���^�����������U�졸�V��H�QV�ҡ���H$�QDV�ҡ���U�H$�AdRV�Ѓ���^]� ��U�졸�V��H�QV�ҡ���H$�QDV�ҡ���U�H$�ARV�Ѓ���^]� ��U�졸�V��H�QV�ҡ���H$�QDV�ҡ���H$�U�ALVR�Ѓ���^]� �̡��V��H$�QHV�ҡ���H�QV�҃�^�������������U�졸��P$�EPQ�JL�у�]� ����U�졸��P$�R]�����������������U�졸��P$�Rl]����������������̡���P$�Bp����̡���P$�BQ�Ѓ����������������U�졸��P$��VWQ�J�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]� ���U�졸��P$�EPQ�J�у�]� ����U�졸��P$��VWQ�J �E�P�ы���u���B�HV�ы���B$�HDV�ы���B$�HLVW�ы���B$�PH�M�Q�ҡ���H�A�U�R�Ѓ� _��^��]� ���U�졸��P$��VWQ�J$�E�P�ы���u���B�HV�ы���B$�HDV�ы���B$�HLVW�ы���B$�PH�M�Q�ҡ���H�A�U�R�Ѓ� _��^��]� ���U���,VW�E�P�o�������Q$�JP�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�ҡ���H$�AH�U�R�Ћ���Q�J�E�P�у� _��^��]� �����̡���P$�B(Q��Yá���P$�BhQ��Y�U�졸��P$�EPQ�J,�у�]� ����U�졸��P$�EPQ�J0�у�]� ����U�졸��P$��VWQ�Jt�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]� ���U�졸��P$�EPQ�J4�у�]� ����U�졸��P$�EPQ�J8�у�]� ����U�졸��UV��H$�ALVR�Ѓ���^]� ��������������U�졸��H�QV�uV�ҡ���H$�QDV�ҡ���H$�U�ALVR�Ћ���E�Q$�J@PV�у���^]�U�졸��UV��H$�A@RV�Ѓ���^]� ��������������U�졸��P$�EPQ�J<�у�]� ����U�졸��P$�EPQ�J<�у����@]� ���������������U�졸��P$�EP�EPQ�JP�у�]� U�졸��P$�EPQ�JT�у�]� ���̡���H$�QX�����U�졸��H$�A\]�����������������U�졸��P$�EP�EP�EPQ�J`�у�]� �����������̡���H(�������U�졸��H(�AV�u�R�Ѓ��    ^]��������������U�졸��P(�R]����������������̡���P(�B�����U�졸��P(�R]�����������������U�졸��P(�R]�����������������U�졸��P(�R ]�����������������U�졸��P(�E�RjP�EP��]� ��U�졸��P(�E�R$P�EP�EP��]� ����P(�B(����̡���P(�B,����̡���P(�B0�����U�졸��P(�R4]�����������������U�졸��P(�RX]�����������������U�졸��P(�R\]�����������������U�졸��P(�R`]�����������������U�졸��P(�Rd]�����������������U�졸��P(�Rh]�����������������U�졸��P(�Rl]�����������������U�졸��P(�Rx]�����������������U�졸��P(���   ]��������������U�졸��P(�Rt]�����������������U�졸��P(�Rp]�����������������U�졸��P(�BpVW�}W���Ѕ�t:����Q(�Rp�GP���҅�t"����P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U�졸��P(�BtVW�}W���Ѕ�t:����Q(�Rt�GP���҅�t"����P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U�졸��P(�BpSVW�}W���Ѕ���   ����Q(�Rp�GP���҅���   ����P(�Rp�GP���҅�tp����P(�Bp�_S���Ѕ�tY����Q(�Rp�CP���҅�tA����P(�Bp��S���Ѕ�t*�OQ��������t��$W��������t_^�   []� _^3�[]� ���U�졸��P(�BtSVW�}W���Ѕ���   ����Q(�Rt�GP���҅���   ����P(�Rt�GP���҅�tp����P(�Bt�_S���Ѕ�tY����Q(�Rt�CP���҅�tA����P(�Bt��S���Ѕ�t*�O0Q���+�����t��HW��������t_^�   []� _^3�[]� ���U�������E�    �E�    �P(�RhV�E�P���҅���   �E���uG����H�A�U�R�Ћ���Q�E�RP�M�Q�ҡ���H�A�U�R�Ѓ��   ^��]� ����Qhmhj  P���   �Ћ�����E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P������3�^��]� ����E��Q�M�j HP�EQ�JP�эU�R�T������   ^��]� �����U�졸���V��H�A�U�R�Ѓ��M�Q������^��u����B�P�M�Q�҃�3���]� ����H$�E�I�U�RP�ы���B�P�M�Q�҃��   ��]� �U��Q����P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U�졸��P(�R8]�����������������U�졸��P(�R<]�����������������U�졸��P(�R@]�����������������U�졸��P(�RD]�����������������U�졸��P(�RH]�����������������U�졸��P(�E�R|P�EP��]� ����U�졸��P(�RL]�����������������U�졸��P(�E���   P�EP��]� �U�졸��E�P(�BT���$��]� ���U�졸��E�P(�BPQ�$��]� ����̡���H(�Q�����U�졸��H(�AV�u�R�Ѓ��    ^]��������������U�졸��P(���   ]��������������U�졸��H(�A]����������������̡���H,�Q,����̡���P,�B4�����U�졸��H,�A0V�u�R�Ѓ��    ^]�������������̡���P,�B8�����U�졸��P,�R<��VW�E�P�ҋu������H�QV�ҡ���H$�QDV�ҡ���H$�QLVW�ҡ���H$�AH�U�R�Ћ���Q�J�E�P�у�_��^��]� �������U�졸��P,�E�R@��VWP�E�P�ҋu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]� ��̡���H,�j j �҃��������������U�졸��P,�EP�EPQ�J�у�]� U�졸��H,�AV�u�R�Ѓ��    ^]�������������̡���P,�B����̡���P,�B����̡���P,�B����̡���P,�B ����̡���P,�B$����̡���P,�B(�����U�졸��P,�R]�����������������U�졸��P,�R��VW�E�P�ҋu������H�QV�ҡ���H$�QDV�ҡ���H$�QLVW�ҡ���H$�AH�U�R�Ћ���Q�J�E�P�у�_��^��]� �������U�졸��H��D  ]��������������U�졸��H��H  ]��������������U�졸��H��L  ]��������������U�졸��H�I]�����������������U�졸��H�A]�����������������U�졸��H�I]�����������������U�졸��H�A]�����������������U�졸��H�I]�����������������U�졸��H���  ]��������������U�졸��H�A]�����������������U���V�u�E�P���+�������Q$�J�E�P�у���u-����B$�PH�M�Q�ҡ���H�A�U�R�Ѓ�3�^��]Ë���Q�J�E�jP�у���u=�U�R��������u-����H$�AH�U�R�Ћ���Q�J�E�P�у�3�^��]Ë���B�HjV�у���u����B�HV�у����I�������Q$�JH�E�P�ы���B�P�M�Q�҃��   ^��]�����������U�졸��H�A ]�����������������U�졸��H�I(]�����������������U�졸��H��  ]��������������U�졸��H��   ]��������������U�졸��H��  ]��������������U�졸��H��  ]��������������U�졸��H�A$��V�U�WR�Ћ���Q�u���BV�Ћ���Q$�BDV�Ћ���Q$�BLVW�Ћ���Q$�JH�E�P�ы���B�P�M�Q�҃�_��^��]������U�졸��H���  ��V�U�WR�Ћ���Q�u���BV�Ћ���Q$�BDV�Ћ���Q$�BLVW�Ћ���Q$�JH�E�P�ы���B�P�M�Q�҃�_��^��]���U�졸��H���  ]��������������U���<���SVW�E�    ��t�E�P�   �������/����Q�J�E�P�   �ы���B$�PD�M�Q�҃��}ࡸ��H�u�QV�ҡ���H$�QDV�ҡ���H$�QLVW�҃���t)����H$�AH�U�R����Ћ���Q�J�E�P�у���t&����B$�PH�M�Q�ҡ���H�A�U�R�Ѓ�_��^[��]���U�졸��H�U���  ��VWR�E�P�ы���u���B�HV�ы���B$�HDV�ы���B$�HLVW�ы���B$�PH�M�Q�ҡ���H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]����������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]�������������̡���H���   ��U�졸��H���   V�uV�҃��    ^]�������������U�졸��P�]�⡸��P�B����̡���P���   ��U�졸��P�R`]�����������������U�졸��P�Rd]�����������������U�졸��P�Rh]�����������������U�졸��P�Rl]�����������������U�졸��P�Rp]�����������������U�졸��P�Rt]�����������������U�졸��P���   ]��������������U�졸��P��  ]��������������U�졸��P�Rx]�����������������U�졸��P���   ]��������������U�졸��P�R|]�����������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P�EPQ��  �у�]� �U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U��E��t ����R P�B$Q�Ѓ���t	�   ]� 3�]� U�졸��P �E�RLQ�MPQ�҃�]� U��E��u]� ����R P�B(Q�Ѓ��   ]� ������U�졸��P�R]�����������������U�졸��P�R]�����������������U�졸��P�R]�����������������U�졸��P�R]�����������������U�졸��P�R]�����������������U�졸��P�R]�����������������U�졸��P�E�R\P�EP��]� ����U�졸��P�E��  P�EP��]� �U�졸��E�P�B ���$��]� ���U�졸��E�P�B$Q�$��]� �����U�졸��E�P�B(���$��]� ���U�졸��P�R,]�����������������U�졸��P�R0]�����������������U�졸��P�R4]�����������������U�졸��P�R8]�����������������U�졸��P�R<]�����������������U�졸��P�R@]�����������������U�졸��P�RD]�����������������U�졸��P�RH]�����������������U�졸��P�RL]�����������������U�졸��P�RP]�����������������U�졸��P���   ]��������������U�졸��P�RT]�����������������U�졸��P�EPQ��  �у�]� �U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P�RX]����������������̡���P���   ��U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]��������������U�졸��P���   ]�������������̡���P���   ��U�졸��P���   ]�������������̡���P���   �ࡸ��P���   �ࡸ��P���   ��U�졸��H���   ]��������������U�졸��H��   ]��������������U�졸��H�U�E��VWRP���  �U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]������������U�졸��H���  ]��������������U�졸��P(�BPVW�}�Q�]���E�$�Ѕ�tM����G�Q(�]�E�BPQ���$�Ѕ�t,����G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U�졸��P(�BTVW�}����$���Ѕ�tE����G�Q(�BT�����$�Ѕ�t(����G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U�졸��P(�BTVW�}����$���Ѕ�tr����G�Q(�BT�����$�Ѕ�tU����G�Q(�BT�����$�Ѕ�t8�OQ���������t)�W0R��������t��HW��������t_�   ^]� _3�^]� ���U�졸��P(�} �R8����P��]� �U�졸��P�BdS�]VW��j ���Ћ���Qhm�p���   h�  V�Ћ�����E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ���Q(�BHV���Ѕ�t ����Q(�E�R VP���҅�t�   �3��EP�������_��^[]� ������U�졸��U�� V��H$�IWR�E�P�ы�����B�P�M�Q�ҡ���H�A�U�RW�Ћ���Q�J�E�P�у��U�R�����������H�A�U�R�Ѓ�_��^��]� ����������̡���P�BVj j����Ћ�^���������U�졸��P�E�RVj P���ҋ�^]� U�졸��P�E�RVPj����ҋ�^]� ����P�B�����U�졸��P���   Vj ��Mj V�Ћ�^]� �����������U�졸��P�EPQ�J�у�]� ����U�졸��P�EPQ�J�у����@]� ���������������U�졸��P�E�RtP�ҋ�����   P�BX�Ѓ�]� ���U�졸��P�E�Rlh#  P�EP��]� ���������������U�졸��P�E�RlhF  P�EP��]� ���������������U�졸��P�E�RtP�ҋ�����   �M�R`QP�҃�]� ���������������U�졸��P���   ]��������������U�졸��P�E���   P�҅�u]� ������   P�B�Ѓ�]� ��������U���V�u�W�}�������Dz�F�G������D{:�G����$�6� �F��$�]��&� �E���������D{_�   ^��]�_3�^��]���������������������U���VW�M��P����E�}��t-����Q4P�B�Ѓ��M��u����_3�^��]Ë�R(�����H0�QW�҃��M��tԋ�R Q�MQ���ҋ���P�B �M��Ѓ��t����Q0�Jx�E�PW�у��M�����_��^��]�������U�졸��P�B VW�}�����=NIVb��   ��   =TCAbtR=$'  t6=MicM��   ����Q���   j hIicM���ЋWP�B����_^]� ��BW����_�   ^]� ����Q���   j hdiem���ЋWP�B����_^]� =INIb��   �~ u���B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� �A�  _3�^]� =cnys����_3�^]� ������V����m����H0�Vh@��҉F���F    ��^�����V��F��m��t����Q0P�B�Ѓ��F    ^�����̡���P0�A���   P�у����������U�졸��P0�E�I���   PQ�҃�]� �������������̡���I�P0���   Q�Ѓ���������̡���P0�A���   j j j j j j j j j4P�у�(������̡���P0�A���   j j j j j j j j j;P�у�(�������U�졸��P0�E�IPQ���   �у�]� ��������������U����E V��P�M��+�������E�Q�R4Ph8kds�M��ҡ���E     �H0���   �U R�U�E�P�Ej R�UP�ER�UP�FRj2P�ыu ��(�M��������^��]� ��������������̡���I�P0���   Q�Ѓ����������U��V��F��u^]� ����Q0�M ���   j j j j j Q�Mj QjP�ҡ���H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uË���Q0P�B�Ѓ������̋A��u� ����Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5���v0Q�MQP���   R�U�R�Ћu�    �F    ������   j P�BV�Ћ�����   �
�E�P�у�$��^��]� �������U�졸��P0�E�I�RPQ�҃�]� �U��A��t)����Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5���v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5���v0QP���   R�Ѓ�^]� �����������U��Q��u3�]� �E�H� V�5���v0Q�MQPR�V\�҃�^]� ����������U��A��u]� ����Q4�M��  Q�MQP�҃�]� �U��A��u]� ����Q4�M�RhQ�MQP�҃�]� ����U��A��u]� ����Q4�M�RpQ�MQP�҃�]� ����U��A��u]� ����Q4�M��  Q�MQP�҃�]� �U���$VW��htniv�M��9�������P�E�R4Phulav�M��ҡ���P�B4hgnlfhtmrf�M��Ћ���E�Q�R4Phinim�M��ҡ���P�E�R4Phixam�M��ҡ���P�E�R4Phpets�M��ҡ���P�E�R4Phsirt�M��ҋE �}$=  �u�����t.����QP�B4h2nim�M��Ћ���Q�B4Wh2xam�M��ЋU�M�QR�E�P������������   P�B8�Ћ�����   �
���E�P�у��M��X���_��^��]�  ��������������U���$V��htlfv�M�������E����P�B,���$hulav�M��Ћ���E,�Q�R4Phtmrf�M����E����P�B,���$hinim�M����E����Q�B,���$hixam�M����E$����Q�B,���$hpets�M��Ћ���ED�Q�R4Phsirt�M����E0��������������Dzw�E8������Dzm�؋���E@�Q�R4Phdauq�M��ҋM�E�PQ�U�R���-���������   P�B8�Ћ�����   �
���E�P�у��M��������^��]�@ �ء���P�B,���$h2nim�M����E8����Q�B,���$h2xam�M����V���U���$V��hgnrs�M��Z����E����E��E�   �Q���   �E�Pj�M��ҡ�����   ��U�R�ЋM����M����E�   �B���   �M�Qj�M��ҡ�����   ��U�R�ЋU���M�QR�E�P������������   P�B8�Ћ�����   �
���E�P�у��M��������^��]� �U���$V��hmnrs�M��z�������P�E�R4Pj�M��ҋM�E�PQ�U�R������������   P�B8�Ћ�����   �
���E�P�у��M��^�����^��]� �����U��E��$�����VDSSS��P�M����������Q�B �M��Ћ���QjP�B4�M��ЋU�M�QR�E�P�������������   P�B8�Ћ�����   �
���E�P�у��M��������^��]� �����������U���$V��hCITb�M��Z�������P�E�R8PhCITb�M��ҡ���P�E�R4Phsirt�M��ҡ���P�E�R4Phulav�M��ҋM�E�PQ�U�R���<���������   P�B8�Ћ�����   �
���E�P�у��M��	�����^��]� U��E��Vj ��P�M�Q�M�����UPR���)�������H�A�U�R�Ѓ���^��]� ����������U��E,��UPj ���T$�$htemf�E$�� �\$�E�\$�E�\$�E�$R�/���]�( �����������U���E����m������m��m��D{���������E����m������D{����E,��Pj ���T$�U�$hrgdf�E$�� �������\$���\$�\$�E�$R����]�( ���������U��E,��Pj ���T$�U�$htcpf�E$�� ��g�����\$�E���\$�}�\$�E�$R�C���]�( ���������������U��Q��u3�]� �E�E�H� V�5���v0Q�M Q�M���\$�E�$QPR�V(�҃�$^]� ������U��Q��u3�]� �E�H� V�5���v0Q�MQPR�V,�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5���v0Q�MQPR�V,�҃�^]� ����������U��Q��u3�]� �E�H� V�5���v0Q�MQPR�V0�҃�^]� ����������U��SVW���W��t$�E�H�5���^0� �uQVP�C0R�Ѓ���u	_^3�[]� �W��t��E�H� ����[0Q�NQPR�S0�҃���t̋W��tŋE�H� �=���0Q��VP�G0R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5���v0Q�MQ�MQPR�V<�҃�^]� ������U��QV3�W��u3��,�E�H� �5���v0Q�MQPR�V,��3Ƀ�9M���������M�B�P0VQ�M�ҋ�_^]� ����U��AV��u3��"�M�Q�	�5���v0R�URQP�F,�Ѓ�������Q�E�M�R4PQ�M�ҋ�^]� ���������������U��A��V��u3��"�M�Q�	�5���v0R�U�RQP�F0�Ѓ�������E��Q�E�M�R,���$P�ҋ�^��]� �����U�����V���U�V�U��]�W��t$�E�H� �=���0Q�M�QPR�W0�҃���u
_3�^��]� �V��t�E�H� �=���0Q�M�QPR�W0�҃���tˋV��tċE�H� �5���v0Q�M�QPR�V0�҃���t�����P�M�RH�E�PQ�M��_�   ^��]� �����������U��� ��A�U�V�U�W�]���u3��&�M�Q�	�5���v0R�U�R�U�RQP�F<�Ѓ����E�}���t����Q�RH�M�QP���ҋE���t����E��Q���$P�B,����_��^��]� U�졸��P�E���   Vj ��MP�ҋM$�U Q�MR�Uj Q�MR�UQPR������^]�  ����������U�졸���P�E���   V���$��MP���E8�E@�M,�Uj P���\$�E0�$Q�E$�� �\$���E�\$�E�\$�$R�����^]�< ������U�졸���P�E���   V���$��MP����Ej j ���T$���$htemf�E$�� �\$�E�\$�E�\$�$P����^]�$ �����������U�졸���P�E���   V���$��MP���E$�Ej �� �\$���E�\$�E�\$�$P����^]�$ ��������������U�졸���P�E���   V���$��MP����j j ���T$�E�$htcpf�E$�� ��g�������\$�E���\$�}�\$�$P����^]�$ ���������������U�졸���0V��H�A�U�WR�Ћ���Q�M���   ���E�PQ�M�E�P�ҋ�����H�A�U�R�Ћ���Q�J�E�PW�ы���B�P�M�Q�ҋE�U��Pj �M�QR����������H�A�U�R�Ћ���Q�J�E�P�у�_��^��]� U���dV��M���������Q���   P�EP�M�Q�M��P�M������M������j j �E�P�M������MPQ������������B�P�M�Q�҃��M������M�������^��]� �����U���P��EV�]���W�}����t����Q���$P���   �����]������U��UЍE��]؋Q�M���   PQ�E�P���ҋ�M��P�U�H�M�P�U�H�M��P�F�U��u_^��]� �M�E�Q�	�5���v0R�U R���\$�U��E��$RQP�F(�Ѓ�$_^��]� ���������������U���0�E�M���u����H���   �҅�u��]� SVW���[  ��htlfv�MЉu�*����E�}����X�U�����$�|{ �]��G�$�n{ �}�S,�M��$hulav�ҡ���P�B4hmrffhtmrf�M��Ћ}�����M�Y���$�%{ �]��G�$�{ �}�S,�M��$hinim�ҋ}�����M�X���$��z �]��G�$��z �}�S,�M��$hixam���衸��P�B,���$hpets�M��Ћ���Q�B4j hdauq�M��Ћ���Q�B4Vhspff�M��Ћ���E �Q�R4Phsirt�M��ҋM�E�PQ�M��U�R����������   P�B8�Ћ�����   �
���E�P�у��M������_��^[��]� U��E��V���u����H���   �҅�u^��]� ����Y  �E�F��u3��"�M�Q�	�5���v0R�U�RQP�F0�Ѓ����E����m�M������\$�M��$� ��M��P�Q�P�Q�@�A��^��]� ����������U���0���]�V���M�]�P���   �E�PQ�M�E�P�ҋ�P�M��Hj �U�P�E P�M��MQ�M�U��UR�U�E�PQR������^��]� ���������������U�����UV�]���E�P�]��ERP��������Q�M�R@���E�PQ�M�ҋ�^��]� ����������U��A��u]� �M�Q�	V�5���v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� ����Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� ����Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U�졸��P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� ����Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj>P�ҋE���(��]� ������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5���v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M�� �MQ�U�R�M��� ��tm�}��E��tN������   P�BH�ЋM��I����tQ�W�7����[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M�� ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5���v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� ����E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� ����Q0�M�RDQ�MQ�MQP�҃�]� U��A��u]�  ����Q0�M$Q�M Q�M���   Q�MQ�MQ�MQ�MQ�MQP�҃�$]�  ��������̋A��uË���Q0P�BX�Ѓ�������U��A��u]� ����Q0�M�RLQ�MQP�҃�]� ����U��A��u]� ����Q0�M�RP��   �QP�҃�]� ��U��A��u]� ����Q0�M�RPQP�҃�]� ��������U��A��u]� ����Q0�M�RTQ�MQ�MQ�MQP�҃�]� ������������U�졸�V�u�VW���H4�R�ЋE�F    �~�H� ����R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� ����Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I����R0P�EPQ���   �у�]� ������̡���I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u���� ����R0�I�R@V�uVP�EPQ�҃�^]� �����������U�졸��P0�E�I�RdP�EP�EP�EP�EPQ�҃�]� �U�졸��P0�E�I�RpP�EP�EP�EP�EPQ�҃�]� �U��E�P� V�5���v0R�UR�UR�UR�URP�A�NhP�у�^]� ��������U��E� ����R0j j j j j j j P�A���   jP�у�(]� �����������U��E� ����R0j j j j j jj P�A���   jP�у�(]� �����������U��E� ����R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M��?����E�H� ����R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R�k����M��S�����^��]� ����������U��E�P� V�5���v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5���v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5���v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5���v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U�졸��P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U�졸��UVj j j j j R��H0�E�Vj P���   jR�Ћ���Q0�E�N�RtPQ�҃�0^]� ��U�졸��P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡���P0�A���   j j j j j j j j jP�у�(�������U�졸��P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡���P0�A���   j j j j j j j j j(P�у�(�������U�졸��P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U�졸��P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡���P0�A���   j j j j j j j j jP�у�(������̡���P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}�M���t����P���   j j���Љ�u��t����Q���   j j���Љ����Q0�E��H�R`VWQ�҃�_^[��]� �U�졸��P0�E�I���   P�EP�EPQ�҃�]� �����̡���P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V����m����H0�Vh@��҉F3��F�F����m�F   ��^�������V��F��m��t����Q0P�B�Ѓ��F    ^������U��V��F�F    ��tn����Q0j j j j j j j j jP���   �Ћ���Q0�E�MP�E���   Q�MP3�9EQ�N��j ��
PQ�҃�D��t�~ t
�   ^]� 3�^]� �������U��E�A�I��u3�]� ����B0Q�H�у�]� ����U�졸��P�B S�]V�����=ckhc��   ��   =cksate=TCAb��   ����Q���   Wj hdiem���Ћ���BSW���F   �Ѓ~ ��t��t��u3Ƀ���Q���C���_^��[]� �~ tn��B����^[]� �~ tY����Q0�F���   j j j j j j j j j P�у�(��t+�F    ^�   []� =atnit�URS���l���^[]� ^3�[]� ��������������U��V��~ ��   W�}����   �$����E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN����M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W��`  ���F    _^]� ĶҶ������-�<�����U��V��~ �  �E W�}�E����   �$�����]������   �   ���]����A��   �   ���]����A��   �t���]������   �b�E������A��uP��������   �E�E��������u3������A{}�,�E���������E������A�����E������DzU����ء���U�H0�F���   j j j j j j j RjP���E �U(��(R���\$�E�$W�_  ���F    _^]�$ �����&�8�U�n�z���������������U���E �E�Uj���\$�E�\$�E�$PR�w���]�  ���U���E �E�Uj���\$�E�\$�E�$PR�G���]�  ���U���E �E�Uj���\$�E�\$�E�$PR����]�  ��̋�3�� �m�H�H�H�������������VW��3���m9~u����H4�V�R�Ѓ��~�~_^����U�졸��P4�E�I�RtPQ�҃�]� �U��U��t3�A����I0R���   P�ҋ���Q0�M���   QP�҃�]� ����P0�E�I�R|PQ�҃�]� ������̡���P4�A�JP�у������������̡���P4�A�JP�у������������̡���P4�A�JP�у������������̡���P4�A�J|P�у������������̡���P4�A���   P�у����������U�졸��E�P4�E$�I��  P�E P�EP�EP���\$�E�$Q�҃�$]�  ��U�졸��P4�E�I�RP�EP�EP�EPQ�҃�]� �����U�졸��P4�E�I�RP�EP�EP�EPQ�҃�]� �����U�졸��P4�E�I�R PQ�҃�]� �U�졸��P4�E�I�R$PQ�҃�]� �U�졸��P0�E�I���   P�EP�EP�EPQ�҃�]� ��U�졸��P0�E�I���   PQ�҃�]� ��������������U�졸��E�P0�E�I���   ���$P�EPQ�҃�]� �U�졸��P4�E�I���   PQ�҃�]� ��������������U�졸��P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U�졸��P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U�졸��P4�E�I�R(PQ�҃�]� �U�졸��P4�E�I�R,P�EP�EPQ�҃�]� ���������U�졸��P4�E�I�R0P�EPQ�҃�]� ������������̡���P4�A�J4P��Y��������������U���S�]V3�����W�~�E�E��QP���   j���Ћ���E��Q���   j j���Ћ���E�Q0�EP�G�M�Q�J`P�ы���B4�N�PQ�ҋ���Q0�Rhj �M�Q�M�Q�M�Q�M�QP�F�HQ�҃�,�} _^[t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� U�졸��P4�E�I�R8PQ�҃�]� �U�졸��P4�E�I�R<PQ�҃�]� �U�졸��P4�E�I���   P�EPQ�҃�]� ����������U�졸��E�P4�A��  ���$P�у�]� ��������̡���P4�A�J@P�у������������̡���P4�A��  P�у����������U�졸��P4�E�I�RDP�EPQ�҃�]� �������������U�졸��P4�E�I�RHP�EPQ�҃�]� �������������U�졸��P4�E�I�RLP�EPQ�҃�]� �������������U�졸��P4�E�I�RPP�EPQ�҃�]� �������������U�졸�SV�uW�����   �QV�҃�����   ������   �]�QS�҃�S��uA������   �Q@�ҋء�����   �Q@V�ҋ���Q4�JPSP�GP�у�_^[]� ������   �H�у���uD������   �H8S�ы���؋��   �H@V�ы���J4�WSP�AHR�Ѓ�_^[]� h(nh�  ��   ������   �BV�Ѓ�����   ������   �]�BS�Ѓ�S��uC������   �B@�Ћ�����   �؋B8V�Ћ���Q4�JLSP�GP�у�_^[]� ������   �H�у���uD������   �H8S�ы���؋��   �H8V�ы���J4�WSP�ADR�Ѓ�_^[]� h(nh�  �
h(nh�  ����Q��0  �Ѓ�_^[]� �U�졸��P4�E�I��  P�EP�EP�EPQ�҃�]� ��U�졸��P4�E,P�E(P�E$P�E �IP�E�RTP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U�졸��P4�E�I�RXP�EP�EP�EPQ�҃�]� ����̡���P4�A�J`P��Y�������������̡���P4�A�JdP�у�������������U�졸��P4�E�I��   P�EP�EP�EPQ�҃�]� ��U�졸��P4�E�I�R\P�EP�EP�EP�EP�EPQ�҃�]� �������������U�졸��P4�E�I�RhP�EPQ�҃�]� �������������U�졸��P4�E�I��  P�EPQ�҃�]� ����������U�졸��P4�E�I��  P�EPQ�҃�]� ����������U�졸��P4�E�I�RpP�EPQ�҃�]� �������������U���,V��~ ��   ����V�H4�AR�Ѓ} t ����Q0�RlP�F�HQ�҃�^��]� ��hARDb�MԉE��E�    輾��P�M�Q�N�U�R�����������   ��U�R�Ѓ��M��;��^��]� ������U�졸��P4�E�I�RlPQ�҃��   ]� ������������U�졸��E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U�졸��P4�E�I���   P�EP�EPQ�҃�]� �����̡���P4�A���   P�у���������̡���P4�A��  P�у���������̸   ����������̸   �����������U�졸�V��H4�V�A$h�  R�Ћ���Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U�졸��P4�E�I�RxP�EP�EP�EPQ�҃�]� �����U�졸��P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}�M���t����P���   j j���Љ�u��t����Q���   j j���Љ����Q4�E��H�RpVWQ�҃�_^[��]� �U��Q����P�B SVW�}���3���=INIb�/  �  =SACbvt+=$'  t
=MicM�  ��B$W����_�   ^��[��]� ��R3��E��E�EP�M�Q���҅�t����U�H4�E�R�VP�AR�Ѓ�_�   ^��[��]� =ARDb�  ����Q���   j j���Ћ���Qj �؋��   j���Ћ���Qj �E����   j���Ћ���Qj �E���   j���ЋM���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>���Y���P���1���P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� ����Q���   j hIicM���ЋWP�B ����_^[��]� �������������U�졸��P4�E�I�RTh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M��z�������Q4�JlP�FP�у��M�蜹��^��]��������V����m����H0�Vh@��҉F���F    �ln�F   ��^��������V��F��m��t����Q0P�B�Ѓ��F    ^������U�졸��P�B VW�}�����=cksat`=ckhct�MQW���ݻ��_^]� �Nj j j j j j �F   ����B0���   j j j Q�҃�(��t'_�F    �   ^]� �~ t��P����_^]� _3�^]� ���U�졸��H���  ]��������������U�졸��H0���   ]��������������U�졸��H0�U�E��VWRP���   �U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]������������U�졸��H0���   ]��������������U�졸��H0���   ]��������������U�졸��H0���   ]��������������U��Ej0P��F  ��]��������������U��Ej0P��  ��P�F  ��]�����U��E�M��j0PQ�U�R��  ��P�nF  ����H�A�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P���  ��P�*F  ����Q�J�E�P�у���]��U��Ej$P�F  3Ƀ�������]����U��Ej$P���  ��P��E  3Ƀ�������]�����������U��E�M��Vj$PQ�U�R���  ��P�E  ���3Ƀ��B�P����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P���  ��P�IE  ���3Ƀ��B�P����M�Q�҃���^��]����U�졸��H�U�E���   RPj �у�]���������������U�졸��H�U�ER�UP���   Rj �Ѓ�]�����������U�졸��P4�E�I�R,P�EP�EPQ�҃�]� ���������U�졸��P4�E�I�R0P�EPQ�҃�]� ������������̡���P4�A�J4P��Y��������������U�������P���   VW�}j ��j���Ћ���E��Q���   j j���Ћ���E�Q0�EP�F�M�Q�J`P�ы���J0�E�P� R�U�R�U�R�U�R�U�R�VP�AhR�Ѓ�(�} _^t&�} t&�E��M�;�~8M�;�}1�E�M�;�~'M���} u�E��M�;�~M�;�}�   ��]� 3���]� ���������������U��ESVW�؅�u�Y����P�}���   j hdiuM���Ћ���tK;3u	_^3�[]� ����Q���   j hIicM����;�u����Q���   j h1icM���Шu��3_^�   []� �����U�졸��P�BT��(V�uhfnic���Ѕ�t����Q�ȋ��   j
�Ѕ���   ����Q�RPhfnic�E�P����P�M��߲���M�������u�E�P��������M���������Q�B ���Ѓ��t����Q�B ���Ѕ�u����Q�B$hfnic���Ћ���E�Q�R8Pj
����^��]���������U�졸��P0�E�IP�EP�EP�EPQ���   �у�]� ��U�졸��P0�E�IV�p� ���   V�uj j j V�uVj Pj=Q�҃�(^]� ����U�졸��P0�E�IV�p� ���   V�uV�uj j j�Vj Pj=Q�҃�(^]� ���̡���I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V����m����H0�WVh@��ҋ}�F�E�F    �F   ��n�F����Q���   ��j hmyal���ЉF��t��t�F    ����Q���   j
hhfed���ЉF_��^]� �����������U�졸��P�B VW�}�����=ytsdt�MQW������_^]� ����B0�N���   Q�ҋ�P������_�   ^]� ��3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ��������������������̸�n�����������U���E�Y(]� ���U���(V���P(�M�Q���ҋN��t&����R0j j j j j j P���   j jQ�Ѓ�(����Q�J�E�P�ы���B�P�M�Q�ҋF����t'����Q0���   j j j �M�Qj jj?j P�҃�$����H�A�U�WR�Ћ���Q�J�E�P�ыF����u3��;����E�    �J0�U�Rj j j h  
 j�U�Rh�  jP���   �Ћ}���(����Q�J�E�P�у���_u3�^��]Ë���B�P�M�Q�ҋF����t'����Q0���   j j j �M�Qj j j8j P�҃�$����H�A�U�R�ЋF����t����Q0jP�BP�Ѓ�����Q�J�E�P�у��M�蛭��Ph   h  K j;�U�Rh	��h�  ���y�������H�A�U�R�Ѓ��M�轭���F��t����Q0P�BX�Ѓ��F��t����Q0P�BX�Ѓ��F��t'����Q0j j j j j jj j jP���   �Ѓ�(j�v$�3<  ���   ^��]�������U���SVW��j�N��  ��V�^(3ۉ^4�^8�^<����H0�Ah�   R�Ћ���Q�J�E�P�ы���B�PSj��M�h�nQ�҃�SS�E�P�M�Q���E��  �]���������B�P�M�Q�҃�Sj�N�K�  _^[��]����̍A�������������U��VW��~4 tA�I ����H��0  h(nh~  ��j
�OE  ����HP�V �AR�Ѓ���uP9F4u���QP�Bh�N0�Ѓ~4 t<����Q��0  h(nh�  �Ћ���QP�Bl���N0���n���_3�^]� �M�U�N8�V4����PP�Bl�N0�Ѓ~4 t%j
�D  ����QP�F �JP�у���u�9F4uۋ���BP�PhS�N0�ҋ^<�F<    ����PP�Bl�N0�Ћ�[_^]� ���U�졸��P�B ��@VW�}�����=MicMtg=ckhctI=fnic��   j�M������uP���&����M���������Q�B4jj����_�   ^��]� ��B�������_��^��]� ����Q���   j hIicM����=�����   htats�M��d�������Q�B0j j�M��ЍM�Q�U�R�E�P���E��  �E�    �n���������   �
�E�P�у��M��O����F�F   ��t����J0�QP�҃��EPW������_^��]� �����������U��E��V��t3�^]� j�N���  j��8  �F    �v����t����H0�QV�҃��   ^]� ��������������j����  j�8  ��3�����������U��E3�h�����h  ���P�Ej BR�Uj PR�ղ��]� �U��Q�Q��u3���]� �E�H� V�5��Q�M�Q�E�    �v0PR�V8�ҋ�����t@�E���t9����Q�M�RQP�ҋE�����t����QW��P�B��W蓃����_��^��]� ������U�졸���V��H�A�U�R�ЋU���M�QR���D�������u����H�A�U�R�Ѓ�3�^��]� �M�Q�M腅������B�P�M�Q�҃���^��]� �������U�졸���V��H�A�U�R�ЋU���M�QR��������M����P�R8�E�PQ�M�ҡ���H�A�U�R�Ѓ���^��]� �������������U���V��M��ς���M�E�PQ�������������B�U�@<�M�Q�MR�ЍM�荃����^��]� ����U�졸��P�E���   Vj ��MP��h���h  �j j jj P�EP���ð��^]� ��������������U�졸�V�uW�����   �QV�҃�V��u,������   �Q@�ҋ���Q4�J P�GP�у�_^]� ������   �H�у���u.������   �H8V�ы���J4�WP�A$R�Ѓ�_^]� ����Q��0  h(nh
  �Ѓ�_^]� �����U���4����H�QSVW�}W�ҡ���P�u���   ��3�SS�Ή]�Ћ���QS�E����   j���Ћ�;��L  �d$ �} ~l����Q�J�E�P�ы���B�Pj j��M�h�nQ�ҡ���P�B<�����Ћ���Q�RLj�j��M�QP���ҡ���H�A�U�R�Ѓ�����Q0�E����   VP�M�Q�ҋ���H�A�U�R�Ћ���Q�J�E�PV�ы���B�P�M�Q�ҡ���P�B<�����Ћ���Q�RLj�j��M�QP���ҡ���H�A�U�R�Ћ���Q�u���   �E��j ��
S���Ћ���Q���   �E�j �CP���ҋ����������_^[��]����������������U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj AQj R�UR������^]� ��������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR语��^]� ����������U��E�E43҃8��R�U<R�U(���\$�E,�$R�E �� �\$�E�\$�E�\$�@�E�$P袮��]�8 ��������������U��E�@3҃8��E��Rj ���T$�$htemf�E �� �\$�E�\$�E�\$�$P�G���]�  ���U��E�E 3҃8��R�� �\$�E�\$�E�\$�@�E�$P����]�  ������U��E�@3҃8��E��Rj ���T$�$htcpf�E �� ��g�����\$�E���\$�}�\$�$P諭��]�  �������U��E3҃8��R�UR�UR�UR�UP�EPR����]� U��E3҃8V�u��V��RP�EP�߰��^]� ����������U��Q��u3�]� �E�E�H� V�5���v0Q�M Q�M���\$���E�$QPR�V(�҃�$^]� ���U�졸��P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U�졸��P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U�졸���P�E���   V���$��MP�ҋ���u�^�    ^]� ��u�F������D{�   ^]� ��^]� ����U���0���U�V�U���M�]��P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�Q�P�Q�P�@�Q�A���O	  ^��]� ��������U���0���]�S��V�]�W��P�M���   �E�PQ�M�E�P�ҋ�x�X��@�U��}�]��E����u�V�~�^_�    �F^[��]� ��u�E�P�NQ��������t�   _^[��]� ������������U���VW�}�M�;}us����P�u���   j htsem���Ѕ�uS����QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E�藰����t�E�M�P�  _�   ^��]� _3�^��]� U��SVW�}��;}u~����P�u���   j htsem���Ѕ�u^����QP���   hrdem���Ѕ�uA�M�E�A��t4����J0j �URWP�A,�Ѓ���t�MQ���  _^�   []� _^3�[]� ���������U���SVW�}��;}��   ����P�u���   j htsem���Ѕ�ug����QP���   hrdem���Ѕ�uJ�M��A�]���t;����J0j �U�RWP�A0�Ѓ���t�E������$�  _^�   [��]� _^3�[��]� �������U���4�ESW�}�M�;�t;Et	;E��   ����P�]���   j htsem���Ѕ���   ����QP���   hrdem���Ѕ�uj�M��U�ỦE��UԉE��]܉E�M�E�P�M�Q�M�U�U�R�E�P�}��Q�����t+�E̋M�������E��X�E��X��  �   _[��]� _3�[��]� ��������U���SVW�}��;}��   ����P�u���   j htsem���Ѕ�uj����QP���   hrdem���Ѕ�uM��U�M��]���Q�M�]��E�R�E�P�}�������t%�E��������E��X�  �   _^[��]� _^3�[��]� ���̋A���X(Q�ȋB$��j j h����.  ���������������U�졸���@VW���H�A�U�R�Ћ���Q�J�E�P�ы���B�U���M�QR���   �M�Q�M�ҋ���H�A�U�R�Ћ���Q�J�E�PV�ы���B�P�M�Q�ҡ���H�I�U�R�E�P�ы���B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�B����V�Ћ���Q�JV�E�P�у����  ����B�P�M�Q�҃�_^��]� ��U���SVW�}��;}��   ����P�u���   j htsem���Ѕ�ue����QP���   hrdem���Ѕ�uH����Q�J�E�P�ыM���U�R�E�P�}��E�    ������u ����Q�J�E�P�у�3�_^[��]� ����B�H����V�ы���B�P�M�VQ�҃����  ����H�A�U�R�Ѓ�_^�   [��]� ������U���V�u3ɍF��H���������M��M����   �RQ�M�QP�ҡ�����   ��U�R�Ѓ���^��]� ����������U���\���SV��H�A�U�WR�Ћ���Q�J3�Sj��E�h oP���F(��g�E��  �]�� 0 ����JP�A(�U�R�Ћ���Q�J���E�P�ы���B�P�M�QW�ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�@�M�Q�U�R�Ћ���Q�B<��8�M��Ћ���Q�RLj�j��M�QP�M���SS�E�P�M�Q���^�������B�P�M�Q�ҡ���H�A�U�R�Ћ���Q�J�E�P�у�htats�M�艘������B�P0jj�M����F(����P�B,���$j�M��ЍM�Q�U�R�E�P���E��  �]��|���������   �
�E�P�у�9^4t[����BP�Ph�N0�ҋF4;�t�N8Q�Ѓ��F<�^8�^4�����B��0  h(nh�  �у�����BP�Pl�N0�ҍM������_^[��]� ����U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�A�E������D{�   ]� ���������U�����u�E�    �Y�E�Y�E�Y]� ��u3�A�E������Dz�A�E������Dz�A�E������D{�   ]� ���������������U��V�����u#�E�M�U�F�E�N�V�    �F^]� ��u�MQ�VR菘������t�   ^]� �������������U��V��F��m��t����Q0P�B�Ѓ��E�F    t	V�(q������^]� ��������������U��V��~ ��mu����H4�V�R�Ѓ��E�F    �F    t	V��p������^]� �������U��V�����u �    ����H�A���UVR�Ѓ��#��u����Q�Rx�EP�N�҅�t�   ����H�A�UR�Ѓ�^]� ������̡���HL���   ��U�졸��H@�AV�u�R�Ѓ��    ^]�������������̡���HL�������U�졸��H@�AV�u�R�Ѓ��    ^]�������������̡���PL���   Q�Ѓ�������������U�졸��PL�EP�EPQ���   �у�]� �������������U�졸�V��HL���   V�҃���u����U�HL���   j RV�Ѓ�^]� ������   �ȋBP�Ћ�����   �MP�BH��^]� �����̡���PL��(  Q�Ѓ�������������U�졸��PL�EP�EPQ��,  �у�]� ������������̡���HL�Q�����U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��PL�E�R��VPQ�M�Q�ҋu��P��腓���M�蝓����^��]� ����U�졸��PL�EPQ���   �у�]� �U�졸��PL�EP�EPQ�J�у�]� ����PL�BQ�Ѓ���������������̡���PL�BQ�Ѓ���������������̡���PL�BQ�Ѓ����������������U�졸��PL�EP�EP�EPQ�J �у�]� ������������U�졸��PL�EPQ��4  �у�]� �U�졸��PL�EP�EP�EPQ�J$�у�]� ������������U�졸��PL�EP�EP�EP�EPQ�J(�у�]� �������̡���PL�B,Q�Ѓ���������������̡���PL�B0Q�Ѓ����������������U�졸��PL�EP�EPQ��  �у�]� ������������̡���PL���   Q�Ѓ�������������U�졸��PL�E��  ��VPQ�M�Q�ҋu��P���b����M��z�����^��]� ̡���PL�B4Q�Ѓ���������������̡���PL�B8j Q�Ѓ��������������U�졸��PL���   ]��������������U�졸��PL���   ]��������������U�졸��PL���   ]��������������U�졸��PL���   ]��������������U�졸��PL���   ]��������������U�졸��PL���   ]��������������U�졸��PL��l  ]��������������U�졸��PL���   ]��������������U�졸��PL���   ]��������������U�졸��PL���   ]��������������U�졸��PL�EPQ�J<�у�]� ���̡���PL�BQ��Y�U�졸��PL�EP�EPQ�J@�у�]� U�졸��PL�Ej PQ�JD�у�]� ��U�졸��PL�Ej PQ�JH�у�]� ��U�졸��PL�EjPQ�JD�у�]� ��U�졸��PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��G  W�M�Q�U�R���$P  ���M����9  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  ��F  j�M�Q�U�R���O  �M���8  ������   ��U�R�Ѓ�^��]�����������U���$����UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��jF  j�E�P�M�Q���	O  �M��a8  ������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}���E  j�E�P�M�Q���N  �M���7  ������   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��E  W�M�Q�U�R���N  ���M����w7  ��t+�u���g��������   ��U�R�Ѓ�_��^[��]� ������   �JL�E�P�ыu��P���h��������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}���D  W�M�Q�U�R���DM  ���M����6  ��t+�u����f��������   ��U�R�Ѓ�_��^[��]� ������   �JL�E�P�ыu��P���Ug��������   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��D  W�M�Q�U�R���L  ���M�����5  _^��[t������   ��U�R�������]Ë�����   �J<�E�P���]�������   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��TC  W�M�Q�U�R����K  ���M����G5  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��B  W�M�Q�U�R���$K  ���M����4  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� �����̡���PL���   Q��Y��������������U�졸��PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U�졸��PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��A  W�M�Q�U�R���I  ���M����3  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��D@  W�M�Q�U�R����H  ���M����72  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��t?  W�M�Q�U�R����G  ���M����g1  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��>  W�M�Q�U�R���$G  ���M����0  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  ��=  j�M�Q�UR���F  �M��/  ������   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��=  j�U�R�E�P���F  �M��v/  ������   �
�E�P�у�^��]� ��������U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���<  j�E�P�M�Q���E  �M���.  ������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��z<  j�E�P�M�Q���E  �M��q.  ������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���;  j�E�P�M�Q���D  �M���-  ������   ��M�Q�҃�_^��]� ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��z;  j�E�P�M�Q���D  �M��q-  ������   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��;  j�U�R�E�P���C  �M��-  ������   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}��:  W�M�Q�U�R���$C  ���M����,  ��t-��u�������   ���^�U�R�Ѓ�_��^[��]� ������   �JP�E�P�ы�u�H��P�@�N����V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���9  W�M�Q�U�R���TB  ���M�����+  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��$9  W�M�Q�U�R���A  ���M����+  ��t������   ��U�R�Ѓ�_^3�[��]Ë�����   �J8�E�P�ы�������   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ���̡���PL���  ��U���$����UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��*8  j�E�P�M�Q����@  �M��!*  ������   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��7  j�U�R�E�P���^@  �M��)  ������   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��O7  h�   �U�R�E�P����?  �M��C)  ������   �
�E�P�у�^��]� �����U�졸��H���   ]��������������U�졸��H���   ]�������������̡���H���   �⡸��H���   ��U�졸��H���   V�u�R�Ѓ��    ^]�����������U�졸��H���   ]��������������U�졸��HL�QV�ҋ���u^]á���H�U�Ej R�UP��h  RV�Ѓ���u����Q@�BV�Ѓ�3���^]��������U�졸��H�U�E��h  j R�U�� P�ERP�у�]����U�졸��H���   ]��������������U�졸��H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡���PL�BLQ�Ѓ���������������̡���PL�BPQ�Ѓ����������������U�졸��PL�EP�EP�EPQ���  �у�]� ���������U�졸��PL�EPQ��  �у�]� �U�졸��PL�EPQ���   �у�]� ̡���PL�BXQ�Ѓ����������������U�졸��PL�EP�EP�EPQ�J\�у�]� ������������U���4���SV��HL�QW�ҋ�3ۉ}�;��x  �M��1{������E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ�����   �BSSW���Ѕ���   ����QL�BW�Ћ���;���   ��    ������   �B(���ЍM�Qh�   ���u��j  ������   �M�;���   ������   ���   S��;�tm������   �ȋB<V�Ћ�����   ���   �E�P�у�;�t����B@�HV�у���;��\����}��M��#  �M��iz����_^[��]� �}�����B@�HW�ы�����   ���   �M�Q�҃��M���"  �M��!z��_^3�[��]� �����̡���PL�B`Q�Ѓ���������������̡���PL�BdQ�Ѓ����������������U�졸��PL�EPQ�Jh�у�]� ���̡���PL��D  Q�Ѓ������������̡���PL�BlQ�Ѓ����������������U�졸��PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh h�
h�
h�
R�Q�U R�UR�UR�U���A�$�5���vLRP���   Q�Ѓ�4^]�  ������̡���PL���   Q�Ѓ�������������U�졸��PL�EP�EP�EPQ��   �у�]� ���������U�졸��PL��H  ]�������������̡���PL��L  ��U�졸��PL��P  ]��������������U�졸��PL��T  ]��������������U�졸��PL��p  ]��������������U�졸��PL��t  ]��������������U�졸��PL�EP�EP�EP�EP�EPQ���   �у�]� �U�졸��PL�EP�EP�EPQ���   �у�]� ���������U�졸��PL�EP�EP�EP�EPQ��   �у�]� �����U�졸��HL���   ]��������������U�졸��HL���   ]��������������U�졸��HL���   ]�������������̡���HL��  �⡸��HL��@  ��U�졸��PL���  ]��������������U�졸��PL���  ]��������������U�졸��PL���  ]��������������U��� ���V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\����QLjP���   ���ЋM��U�Rh=���M�}��  ��������   ���   �U�R�Ѓ��M��u��  ��_^��]Ë�����   ���   �E�P�у��M��u���  _�   ^��]����U��� ���V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\����QLjP���   ���ЋM��U�Rh<���M�}��C  ��������   ���   �U�R�Ѓ��M��u��L  ��_^��]Ë�����   ���   �E�P�у��M��u��  _�   ^��]����U�졸��P8�EPQ�JD�у�]� ���̡���H8�Q<�����U�졸��H8�A@V�u�R�Ѓ��    ^]�������������̡���H8�������U�졸��H8�AV�u�R�Ѓ��    ^]��������������U�졸��P8�EP�EP�EPQ�J�у�]� ������������U�졸��P8�EP�EPQ�J�у�]� ����P8�BQ�Ѓ����������������U�졸��P8�EPQ�J �у�]� ����U�졸��P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U�졸��P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U�졸��P8�EP�EPQ�J(�у�]� U�졸��P8�EP�EP�EPQ�J,�у�]� ������������U�졸��P8�EP�EP�EPQ�J�у�]� ������������U�졸��P8�EP�EP�EP�EP�EPQ�J�у�]� ����U�졸��P8�EP�EPQ�J0�у�]� U�졸��P8�EP�EP�EPQ�J4�у�]� ������������U�졸��P8�EPQ�J8�у�]� ����U�졸��H��x  ]��������������U�졸��H��|  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H�A,]�����������������U�졸��H���  ]��������������U�졸��H�QV�uV�ҡ���H�Q8V�҃���^]�����̡���H�Q<�����U�졸��H�I@]����������������̡���H�QD����̡���H�QH�����U�졸��H�AL]�����������������U�졸��H�IP]�����������������U�졸��H��<  ]��������������U�졸��H��,  ]��������������U�졸��H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡���H���   �⡸��H���  ��U�졸��H�U�ER�UP�ER�UP���   Rh�6  �Ѓ�]����������������U�졸��H�A]�����������������U�졸��H��\  ]��������������U�졸��H�AT]�����������������U�졸��H�AX]�����������������U�졸��H�A\]����������������̡���H�Q`�����U�졸��H���  ]�������������̡���H�Qd����̡���H�Qh�����U�졸��H�Al]�����������������U�졸��H�Ap]�����������������U�졸��H�At]�����������������U�졸��H��D  ]��������������U�졸��H��  ]��������������U�졸��H�Ix]�����������������U�졸��H��@  ]��������������U��V�u���bH������H�U�A|VR�Ѓ���^]���������U�졸��H���   ]��������������U�졸��H��h  ]��������������U�졸��H��d  ]��������������U�졸��H���  ]�������������̡���H���   ��U�졸��H��l  ]��������������U�졸��H��   ]��������������U�졸��H��  ]��������������U��V�u����k������H���   V�҃���^]���������̡���H��`  ��U�졸��H��  ]��������������U�졸��H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U�졸��H���  ]��������������U��U�E����H�E���   R���\$�E�$P�у�]�U�졸��H���   ]��������������U�졸��H���   ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���   ]��������������U�졸��H���   ]��������������U�졸��H���   ]��������������U�졸��H���   ]��������������U�졸��H���   ]��������������U�졸��H���   ]��������������U�������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�������P�E�P�E�P�E�PQ���   �у����#E���]����������������U�졸��H��8  ]��������������U��V�u(V�u$�E�@����R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@����R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U�졸��P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U�졸��P0�EP�EP�EP�EPQ���   �у�]� ����̡���P0���   Q�Ѓ�������������U�졸��P0�EP�EPQ���   �у�]� �������������U�졸��P0�EP�EP�EP�EPQ���   �у�]� ����̡���P0���   Q�Ѓ������������̡���H0���   ��U�졸��H0���   V�u�R�Ѓ��    ^]�����������U�졸��H��H  ]��������������U�졸��H��T  ]�������������̡���H��p  �⡸��H���  ��U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H�U�E��X  ��VR�UPR�E�P�ыu�    �F    ������   �Qj PV�ҡ�����   ��U�R�Ѓ� ��^��]��������U���4VhLGOg�M��\e������Q��X  3�VP�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�у� �M��Be��������   �PT�M�Q�҃���u'�u���d��������   ��U�R�Ѓ���^��]Ë�����   �JT�E�P�ыu��P���d��������   ��M�Q�҃���^��]���������������U�졸��H��  ]��������������U�졸��H��\  ]��������������U�졸��H�U��t  ��V�uVR�E�P�у�����@���M��+@����^��]�����U�졸��H�U���  ��VWR�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]����������������U�졸��H�U���  ��VWR�E�P�ы���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]����������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H�U�E��VWj R�UP�ERP��t  �U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�(_��^��]��U�졸��H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    ������   j P�BV�Ћ�����   �
�E�P�у�$��^��]���U�졸��H��8  ]��������������U���  ���3ŉE��M�EPQ������h   R�`� ����x	=�  |#�����H��0  h0ohH  �҃��E� ����H��4  ������Rhto�ЋM�3̓��t�  ��]�������U�졸��H��  ��V�U�WR�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]����U�졸��H��  ��V�U�WR�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]����U�졸��H��p  ��4�҅���   h���M���_������P�E�R4Ph���M��ҡ���P�E�R4Ph���M��ҡ���H��X  j �U�R�E�hicMCP�ы���E�    �E�    ���   j P�A�U�R�Ћ�����   �
�E�P�ы�����   ��M�Q�҃�$�M��_����]��������U�졸��H��p  ��4V�҅�u����H�u�QV�҃���^��]�Wh!���M���^������P�E�R4Ph!���M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �PH�M�Q�ҋu������H�QV�ҡ���H�QVW�ҡ�����   ��U�R�Ѓ�4�M��}^��_��^��]������U�졸��H��p  ��4V�҅�u����H�u�QV�҃���^��]�Wh����M���]������P�E�R4Ph����M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �PH�M�Q�ҋu������H�QV�ҡ���H�QVW�ҡ�����   ��U�R�Ѓ�4�M��m]��_��^��]������U�졸��H��p  ��4�҅�u��]�Vh#���M���\������P�E�R4Ph#���M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �P8�M�Q�ҋ�����   ��U�R�Ѓ�(�M��\����^��]���������������U�졸��H��p  ��4�҅�u��]�Vhs���M��\������P�E�R4Phs���M��ҡ���H��X  3�V�U�R�E�hicMCP�ы���u��u����   VP�A�U�R�Ћ�����   �
�E�P�ы�����   �P8�M�Q�ҋ�����   ��U�R�Ѓ�(�M��[����^��]���������������U�졸��H���  ]��������������U�졸��H��@  ]��������������U�졸��H���  ]��������������U��V�u���t����QP��D  �Ѓ��    ^]������U�졸��H��H  ]��������������U�졸��H��L  ]��������������U�졸��H��P  ]��������������U�졸��H��T  ]��������������U�졸��H��X  ]��������������U�졸��H��\  ]�������������̡���H��d  ��U�졸��H��h  ]��������������U�졸��H��l  ]�������������̡���H���  ��U�졸��H�U���  ��VR�E�P�ыu��P���Y���M��Y����^��]�����U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H��l  ]��������������U�졸��H���  ]��������������U�졸��H���  ]��������������U�졸��H��$  ]��������������U�졸��H��(  ]��������������U�졸��H��,  ]�������������̡���H��0  �⡸��H��<  ��U�졸��H���  ]�������������̡���H���  ��U�졸��H���  ]������������������������������U�졸��H��  ]�������������̡���H��P  ��U�졸��H��`  ]�������������̡�����   ���   ��Q��Y��������U�졸��H�A�U��� R�Ћ���Q�Jj j��E�hxoP�ы���B�P�M�Q�ҡ���H�I�U�R�E�P�ы���B�P<�� �M��ҋ���Q�M�RLj�j�QP�M��ҡ���H�A�U�R�Ћ���Q�J�E�P�ы���B�P�M�Q�҃���]��������������h��PhD 萅  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h��jhD 輄  ����t
�@��t]��3�]��������Vh��j\hD ��茄  ����t�@\��tV�Ѓ���^�����Vh��j`hD ���\�  ����t�@`��tV�Ѓ�^�������U��Vh��jdhD ���)�  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh��jhhD ����  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh��jlhD ��謃  ����t�@l��tV�Ѓ�^�������U��Vh��h�   hD ���v�  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh��h�   hD ���&�  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh��jphD ���ق  ����t�@p��t�MQV�Ѓ�^]� ���^]� ��U��Vh��jxhD ��虂  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh��j|hD ���Y�  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh��j|hD ����  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� �������������U���Vh��h�   hD ���Á  ����t=���   ��t3�MQ�U�VR��h��j`hD 薁  ����t�@`��t	�M�Q�Ѓ���^��]� �����̋���������������h��jhD �O�  ����t	�@��t��3��������������U��V�u�> t+h��jhD ��  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h��jhD �р  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh��jhD ��艀  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh��jhD ���I�  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh��j hD ����  ����t�@ ��tV�Ѓ�^�3�^���Vh��j$hD ����  ����t�@$��tV�Ѓ�^�3�^���U��Vh��j(hD ���  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh��j,hD ���Y  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh��j(hD ���  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh��j4hD ����~  ����t�@4��tV�Ѓ�^�3�^���U��Vh��j8hD ���~  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh��j<hD ���I~  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh��jDhD ���~  ����t�@D��tV�Ѓ�^�3�^���U��Vh��jHhD ����}  ����t�M�PHQV�҃�^]� U��Vh��jLhD ���}  ����u^]� �M�PLQV�҃�^]� �����������U��Vh��jPhD ���i}  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh��jThD ���,}  ����u^Ë@TV�Ѓ�^���������U��Vh��jXhD ����|  ����t�M�PXQV�҃�^]� U��Vh��h�   hD ����|  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh��h�   hD ���v|  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh��h�   hD ���&|  ����u^]� �M���   QV�҃�^]� �����U��Vh��h�   hD ����{  ����u^]� �M���   QV�҃�^]� �����U��Vh��h�   hD ���{  ����u^]� �M���   QV�҃�^]� �����U��Vh��h�   hD ���f{  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh��h�   hD �%{  ����u����H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ���Q�u���BV�Ћ���Q�BVW�Ћ���Q�J�E�P�у�_��^��]��U��Vh��h�   hD ���z  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   hD ���Fz  ����t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   hD ���z  ����t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   hD ����y  ����t���   ��t�MQ����^]� 3�^]� �Vh��h�   hD ���y  ����t���   ��t��^��3�^����������������U��Vh��h�   hD ���Fy  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh��h�   hD ����x  ����t���   ��t�MQ����^]� ��������U��Vh��h�   hD ���x  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh��h�   hD ���ix  ����t���   ��t��^��3�^����������������VW��3����$    �h��jphD �x  ����t�@p��t	VW�Ѓ������8 tF��_��^�������U��SW��3�V��    h��jphD ��w  ����t�@p��t	WS�Ѓ������8 tqh��jphD �w  ����t�@p��t�MWQ�Ѓ�������h��jphD �kw  ����t�@p��t	WS�Ѓ�����V���������tG�]����E^��t�8��~=h��jphD �w  ����t�@p��t	WS�Ѓ������8 u_�   []� _3�[]� ����������U��Vh��j\hD ����v  ����t3�@\��t,V��h��jxhD �v  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh��j\hD ���iv  ����t3�@\��t,V��h��jdhD �Gv  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh��j\hD ���v  ����tG�@\��t@V�ЋEh��jdhD �E��E�    �E�    ��u  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh��j\hD ���u  ����t\�@\��tUV��h��jdhD �gu  ����t�@d��t
�MQV�Ѓ�h��jhhD �>u  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh��j\hD ����t  ������   �@\��t~V��h��jdhD ��t  ����t�@d��t
�MQV�Ѓ�h��jhhD �t  ����t�@h��t
�URV�Ѓ�h��jhhD �t  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh��jthD ���Ft  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h��j`hD �t  ����th�@`��ta�M�Q�Ѓ���^��]� h��j\hD ��s  �u����t4�@\��t-V��h��jdhD �s  ����t�@d��th��V�Ѓ���^��]� ������U���Vh��h�   hD �us  ����tU���   ��tK�M�UQR�M�Q�Ћu��P���h���h��j`hD �7s  ����te�@`��t^�U�R�Ѓ���^��]�h��j\hD �s  �u����t3�@\��t,V��h��jxhD ��r  ����t�@x��t
�MVQ�Ѓ���^��]�����U���Vh��h�   hD ���r  ����tR���   ��tH�MQ�U�R���ЋuP������h��j`hD �jr  ����t|�@`��tu�M�Q�Ѓ���^��]� h��j\hD �E�    �E�    �E�    �$r  �u����t3�@\��t,V��h��jdhD ��q  ����t�@d��t
�U�RV�Ѓ���^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t������   P�B@��]� �E��t������   P�BD��]� ������   R�PD��]� �����U�졸��P@�Rd]�����������������U�졸��P@�Rh]�����������������U�졸��P@�Rl]�����������������U�졸��P@���   ]��������������U�졸����   ���   ]�����������U�졸����   ���   ]����������̡���P@�Bt����̡���P@�Bx�����U�졸��P@�R|]����������������̡���P@���   �ࡸ����   �Bt��U�졸��P@���   ]�������������̡���P@���   ��U�졸��P@���   ]��������������U�졸��P@���   ]��������������U�졸��P@���   ]��������������U�졸��P@���   ]��������������U�졸��P@���   ]��������������U�졸��P@���   ]��������������U�졸�V��H@�QV�ҋM����t��#�������Q@P�BV�Ѓ�^]� �̡���PH���   Q�Ѓ�������������U�졸��P@�EPQ�JL�у�]� ���̡���P@�BHQ�Ѓ����������������U�졸��P@�EP�EP�EPQ�J�у�]� ������������U�졸��P@�EPQ�J�у�]� ����U�졸��P@�EP�EPQ�J�у�]� U�졸��P@�EPQ�J �у�]� ����U�졸����   �R]��������������U�졸����   �R]��������������U�졸����   �R ]��������������U�졸����   ���   ]�����������U�졸����   ��D  ]�����������U�졸��E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U�졸����   ���   ]����������̡�����   �B$�ࡸ��H@�Q0�����U�졸��H@�A4j�URj �Ѓ�]����U�졸��H@�A4j�URh   @�Ѓ�]�U�졸��H@�U�E�I4RPj �у�]�̡���H|�������U��V�u���t����Q|P�B�Ѓ��    ^]��������̡���H|�Q �����U��V�u���t����Q|P�B(�Ѓ��    ^]��������̡���H@�Q0�����U��V�u���t����Q@P�B�Ѓ��    ^]���������U�졸��H@���   ]��������������U��V�u���t����Q@P�B�Ѓ��    ^]��������̡���PH���   Q�Ѓ�������������U�졸��PH�EPQ��d  �у�]� �U�졸��H �IH]�����������������U��}qF uHV�u��t?������   �BDW�}W���Ћ���Q@�B,W�Ћ���Q�M�Rp��VQ����_^]����������̡���P@�BT�����U�졸��P@�RX]�����������������U�졸��P@�R\]����������������̡���P@�B`�����U�졸��H��T  ]��������������U�졸��H@�U�A,SVWR�Ћ���Q@�J,���EP�ы���Z��h��hE  �΋���;��Ph��hE  ����;��P��T  �Ѓ�_^[]����U�졸��PT�EP�EPQ�J�у�]� U�졸��PT�EPQ�J�у�]� ����U�졸��PT�EPQ�J�у�]� ����U�졸��PT�E�R<��PQ�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�졸��HT�]��U�졸��H@�AV�u�R�Ѓ��    ^]�������������̡���HT�hG  �҃�������������U�졸��H@�AV�u�R�Ѓ��    ^]�������������̡���PD�BQ�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�BQ�Ѓ����������������U�졸��PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U�졸��PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�졸��PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�졸��PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U�졸��PX�EPQ�J�у�]� ����U�졸��PX�EPQ�J�у�]� ����U�졸��PX�EPQ�J�у�]� ����U�졸��PX�EPQ�J�у�]� ����U�졸��PX�EPQ�J$�у�]� ����U�졸��PX�EPQ�J �у�]� ����U�졸��PD�EP�EPQ�J�у�]� U�졸��HD�U�j R�Ѓ�]�������U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��HD�	]��U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��HD�U�j R�Ѓ�]�������U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��U�HD�Rh2  �Ѓ�]����U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��U�HD�RhO  �Ѓ�]����U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��U�HD�Rh'  �Ѓ�]����U�졸��H@�AV�u�R�Ѓ��    ^]�������������̡���HD�j h�  �҃�����������U�졸��H@�AV�u�R�Ѓ��    ^]�������������̡���HD�j h:  �҃�����������U�졸��H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E�������   �R�E�Pj�����#E���]�̡���HD�j h�F �҃�����������U�졸��H@�AV�u�R�Ѓ��    ^]�������������̡���HD�j h�_ �҃�����������U�졸��H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E�����E�    ���   �R�E�Pj������؋�]� ̡���PD�B$Q�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ���������������̡���PD�B(Q�Ѓ���������������̡���PD�BQ�Ѓ����������������U�졸��H �Ah]�����������������U�졸��H@�AV�u�R�Ѓ��    ^]�������������̡���H �������U��V�u���t����Q P�B�Ѓ��    ^]���������U�졸��P �EPQ�J4�у�]� ����U�졸��P �EPQ�J�у�]� ����U�졸��P �EPQ�J�у�]� ���̡���P �BQ��Y�U��V�uW�����/������H �QVW�҃�_��^]� �����U�졸��P �EPQ�J �у�]� ���̡���P �B,Q�Ѓ���������������̡���P �B0Q�Ѓ���������������̡���H\�������U�졸��H\�AV�u�R�Ѓ��    ^]�������������̡���P\�BQ�Ѓ���������������̡���P\�BQ�Ѓ����������������U�졸��P\�EPQ�J�у�]� ����U�졸��P\�EP�EPQ�J�у�]� U�졸��P\�EPQ�J�у�]� ���̡���P\�BQ�Ѓ����������������U�졸��P\�EPQ�J �у�]� ����U�졸��P\�EP�EPQ�J$�у�]� U�졸��P\�EP�EP�EP�EPQ�J`�у�]� ��������U�졸��P\�EPQ�J0�у�]� ����U�졸��P\�EPQ�J@�у�]� ����U�졸��P\�EPQ�JD�у�]� ����U�졸��P\�EPQ�JH�у�]� ���̡���P\�B4Q�Ѓ����������������U�졸��P\�EP�EPQ�J8�у�]� U�졸��P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu��$������H\�QV�҃���S���$��3���~B��I ����H\�U�R�U��EP�A`h���VR�ЋM��Q���c$���U�R���X$��F;�|�_^[��]� ����������U���VW�}�E��P��� ���}� ��   ����Q\�BV�Ѓ��M�Q���a ���E���t]S3ۅ�~H�I �UR���E ���E�P���: ���E;E�!������Q\P�BV�ЋE@���E;E�~�C;]�|�[_�   ^��]� _�   ^��]� U�졸��E�PH�B���$Q�Ѓ�]� ���������������U�졸��PH�EPQ���   �у�]� �U�졸��PH�EPQ���  �у�]� �U�졸��PH�EPQ���  �у�]� �U�졸��PH�EP�EPQ��  �у�]� �������������U�졸��PH�EP�EPQ��  �у�]� ������������̡���PH���  Q�Ѓ�������������U�졸��PH�EPQ���  �у�]� ̡���PH���   j Q�Ѓ�����������U�졸��PH�EPj Q���   �у�]� ��������������̡���PH���   jQ�Ѓ�����������U�졸��PH�EPjQ���   �у�]� ��������������̡���PH���   jQ�Ѓ����������U�졸��PH�EPjQ���   �у�]� ���������������U�졸��PH�EP�EPQ���   �у�]� �������������U�졸��PH�EP�EPQ���   �у�]� ������������̡���PH���   Q�Ѓ�������������U�졸��PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP��� ���������t�E����QH���   PVW�у���_^]� �����U��EVW���MPQ�,���������t�M����BH���   QVW�҃���_^]� ̡���PH���   Q�Ѓ������������̡���PH���   Q�Ѓ�������������U�졸��PH�EPQ���   �у�]� �U�졸��PH�EP�EPQ���  �у�]� �������������U�졸��PH�EPQ���   �у�]� �U�졸��PH�EP�EPQ��8  �у�]� �������������U�졸��PH�EP�EPQ��   �у�]� ������������̡���PH���  Q�Ѓ������������̡���PH���  Q�Ѓ������������̡���PH���  Q�Ѓ������������̡���PH��  Q�Ѓ������������̡���PH��  Q�Ѓ�������������U�졸��PH�EP�EPQ��  �у�]� �������������U�졸��PH�EP�EP�EPQ��   �у�]� ���������U�졸��PH�EP�EP�EP�EPQ��|  �у�]� �����U�졸��PH�EPQ��  �у�]� ̡���PH��T  Q�Ѓ�������������U�졸��PH�EP�EPQ��  �у�]� �������������U�졸��PH�EPQ��8  �у�]� �U�졸��PH�EPQ��<  �у�]� �U�졸��PH�EP�EP�EPQ��@  �у�]� ���������U�졸��PH�EPQ���  �у�]� ̡���PH��L  Q��Y��������������U�졸��PH�EPQ��H  �у�]� ̡��V��H@�Q,WV�ҋ���Q��j �ȋ��   h�  �Ћ���QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡���P@�B,Q�Ћ���Q��j �ȋ��   h�  �������U�졸��E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�졸��E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�졸��PH�EP�EP�EPQ��   �у�]� ��������̡���HH��  ��U�졸��HH��  ]��������������U�졸��E�PH��$  ���$Q�Ѓ�]� �����������̡���PH��(  Q�Ѓ�������������U�졸��PH�EP�EPQ��,  �у�]� �������������U�졸��E�PH�EP�E���$PQ��0  �у�]� ���̡���PH���  Q�Ѓ������������̡���PH��4  Q�Ѓ������������̋��     �������̡���PH���|  jP�у���������U�졸��UV��HH��x  R��3Ƀ������^��]� ��̡���PH���|  j P�у��������̡���PH��P  Q�Ѓ������������̡���PH��T  Q�Ѓ������������̡���PH��X  Q�Ѓ�������������U�졸��PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡���PH��`  Q�Ѓ�������������U�졸��PH�EPQ��d  �у�]� �U�졸��E�PH��h  ���$Q�Ѓ�]� ������������U�졸��E�PH��t  ���$Q�Ѓ�]� ������������U�졸��E�PH��l  ���$Q�Ѓ�]� ������������U�졸��PH�EPQ��p  �у�]� �U�졸��PH�EP�EP�EP�EPQ���  �у�]� �����U�졸��PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U�졸��E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E����HH�E���   R�U���$P�ERP�у�]����������������U���E�M��o輵  �M;�|�M;�~��]�����������U�졸��PH�E���   Q�MPQ�҃�]� ������������̡���PH���   Q��Y�������������̡���PH���   Q�Ѓ������������̡���PH���   Q��Y��������������U�졸��PH�EP�EPQ���   �у�]� �������������U�졸��PH�EP�EP�EP�EP�EPQ���  �у�]� ̡���PH��t  Q��Y�������������̋�� �o�@    ���o����Pl�A�JP��Y��������U�졸�V��Hl�V�AR�ЋE����u
�   ^]� ����Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË���QlP�B�Ѓ�������U�졸��Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E����HH�ER�U���$P���  R�Ѓ�]����U�졸��HH���  ]��������������U�졸��HH���  ]��������������U��U0�E(����HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U�졸��HH���  ]��������������U�졸��E�PH�EP���$Q���  �у�]� ��������U���V�������E����   �} ��   ����HH��p  SWj h�  V�ҋء���HH���   h�  V�]��ҋ������}����   �M3��u���������   �]�E�P�M�Q�MWV�J�����t\�u�;u�T������u�E����ҋL�;L�t-����Bl�S�@����QR�ЋD������t	�M�P�3���F;u�~��}�u�MF�u������;��w����E�_[^��]� 3�^��]� ��������������U������SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u����HH���  �'��u����HH���  ���uš���HH���  S�ҋȃ��E��t�W���������HH���   h�  S3��҃����  ���_�u����    ����Hl�U�B�IWP�ы�������   ����F�J\�UP�A,R�Ѓ���t�K�Q�M���������F�J\�UP�A,R�Ѓ���t�K�Q�M�����E��;Pt&�F����Q\�J,P�EP�у���t	�MS��������v�B\�M�P,VQ�҃���t�M�CP�c�������QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U�졸��HH���   ]�������������̡���PH���   Q��Y��������������U�졸��HH���  ]��������������U�졸���P���   V�uW�}���$V�����E������At���E������z����؋���Q�B,���$V����_^]����������������U���0���U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١���]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U�졸��HH�]��U�졸��H@�AV�u�R�Ѓ��    ^]�������������̡���HH�h�  �҃�������������U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��HH�Vh  �ҋ�������   �EPh�  � �������t]����QHj P���   V�ЋMQh(  ���������t3����JH���   j PV�ҡ�����   �B��j j���Ћ�^]á���H@�QV�҃�3�^]�������U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��HH�Vh�  �ҋ�����u^]á���HH�U�E��  RPV�у���u����B@�HV�у�3���^]�������U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��HH�I]�����������������U�졸��H@�AV�u�R�Ѓ��    ^]��������������U�졸��PH�EPQ���  �у�]� �U�졸��PH�EPQ���  �у�]� ̡���PH���  Q�Ѓ�������������U�졸��HH���  ]��������������U�졸��E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡���PH���  Q�Ѓ�������������U�졸��PH�EP�EPQ���  �у�]� ������������̡���PH��  Q�Ѓ�������������U�졸��PH�EP�EP�EPQ���  �у�]� ��������̡���PH���  Q�Ѓ������������̡���PH���  Q�Ѓ�������������U�졸��PH�EPQ��  �у�]� �U�졸��PH�EPQ��  �у�]� ̋������������������������������̡���HH���  ��U�졸��HH���  ]��������������U�졸��PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U�졸��PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡���PH��,  Q�Ѓ�������������U�졸��PH�EPQ��X  �у�]� ̡���PH��\  Q�Ѓ�������������U�졸��HH��0  ]��������������U�졸���W���HH���   j h�  W�҃��} u�   _��]� Vh�  ������������   ����HH���   j VW�҃��M��������P�E�R0Ph�  �M����E����P�B,���$h�  �M��Ћ���Q@�J(j �E�PV�у��M����^�   _��]� ^3�_��]� �����U��S�]�; VW��u7����U�HH���   RW�Ѓ���u����QH���   jW�Ѓ���t�   �����   ����QH���   W�Ѓ��} u(����E�QH�M���  P�ESQ�MPQW�҃��B�u��t;����U�HH�ER�USP���  VRW�Ћ�����   �B(�����Ћ���uŃ; u����QH���   W�Ѓ���t3���   �W��u1����QH���   �Ћ���E�QH���   PW�у�_^[]� ����BH���   �у��} u0����M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ����QH�h  �Ћ؃���u_^[]� ������   �u�Bx���Ћ�����   P�B|���Ѕ�tU����E�QH�MP�Ej Q���  VPW�у���t������   �ȋBHS�Ћ�����   �B(���Ћ���u�_^��[]� ��������������U��EV���u����HH���  �'��u����HH���  ���u����HH���  V�҃���u3�^]� P�EP���.���^]� ���������U���D����HH���   SV�uWh�  V�ҋء���HH���   3�Wh�  V�]؉}��҉E�3����E�E�E�;���	  ������   �B���Ћ��=�  ��  �QH���   3�Sh:  V�Ћ���QH�E����   h�  V�Ћ���QHS�����   h�  V�}Љ]��Ћ���QH�E䋂  V�Ћ���QH�E̋��  V�Ѓ�(�Eȅ��}   �M���M܋��M̅�tMj�S�L  ���t@�@�Eȃ|� �<�~����%�������;�u/����V  ;E�~�Eԋ��V  E���E܋;Pu�E���E��E�C;]�|��}� t{�}�j V����������  ��������t[���1����]�;�uP����H���  �<[�h�o��h�  W�҃��E���H  �M��E��=���WP�E�P�r�  ����]؋���Q���  �<[�h�o��h�  W�Ѓ��E����  �M�WQP�,�  �E�3ۃ�;�~-����J���   h�o��h�  P�҃��E�;���  ����U�HH��  j�RV�Ѓ�����  �}�;�tjV���������x  �������E���]�����QH���   Sh�  V�Ѓ�3��E��]�9]��Z  �}���}čd$ �M̅��L  �U�j�R�J  ����8  �Mȍ@�|� ���]�~����%�������9E���  ���T  �E�3�3ɉE؉M�9C��   ��$    �����������ti�]������������M�ҋ9�<��}�҉T��y�]��|��]��z�|��y�]��|��]��z�|��I�}��]܉L��M��}ă��T����M�A�M�;K�v����Eԅ��2  �+�����~�M�QPQ�M��	  �U��v�E�3�+M܉E��U�;U���   �}� �E����E�t4M��@�E�Ћ��P�Q�P�Q�P�Q�P�Q�@�A�M܋Eč@�E�Ћ��P�Q�P�Q�P�Q�P�Q�@�A;]�}_�UċE�9�uT�ȋL�����������w0�$�(��U���4���M���t���U���t��	�M���t��M܃�;]�|��E؃�F�M�;]������U�;U��  �U�R������E�P�����M�Q������_^3�[��]Ë�M�3�;G�Å���   �E��v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q�P �Q�P$�Q�P(�I�H,��@�E�ЋU��Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU��Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U�@�ʋU��v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U�@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU��v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U�@�ʋU��v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@���E�}�;E�������U�R�����E�P��������  ���   �B����=  ��  ����QH���   j h(  V�Ћ���QH�؋��   h(  V�ЋЃ�3��Uԅ�~ ��Å�t�|� t�<O��|O�@;�|�}�}؋���Q���  �<�h�o��hY  W�Ѓ��E���   �M�WQP�P�  �}ԋ���B���  �h�o��h^  W�у��E���tEWSP��  �M���+���RH��PQ�E���   V�Ѓ���u�M�Q�x����U�R�o�����_^3�[��]á���HH���   j h�  V�҉E���HH���   j h(  V��3�3���3��Eĉ}��]�9]��8  �U����څ��  �E�    ����   �U��<��v��   ����U�:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U�\�EЉY�\�T�Y�Z�Y �Z�Y$�Z�Y(�R�]�Q,�U�@����0��;�|��}��|� tt�U�M�ύI�ʋU��v���A�B�A�B�A�B�A�B�I�J�E��ЋE��Tv�Ћ��A�B�A�B�A�B�A�B�I�J�U���<ډ}�C�]�;]�������M�3�3�;�~�Uĉt���   @;�|��U�R�������E�P������_^�   [��]ÍI �z�z�z�z��������U��E�MSVW�}�����9|���I ��;|�;�s$���p��Y�X��q;�u����;�uǋ���_^[]� ����������U���W�}����   �Ǚ+���@S�]� �M���V�E��M�\����E��M��I ��~H���m��E��&�s����u�1�3�q�sO��U�M�Q��~S�Ћ�9}���Eҋ�L��;�}�;A}B���;}��E��F�E���A�F�E���E�A�;�~��j���^[_��]� ������������U��V��V��o����Hl�AR�Ѓ��Et	V��������^]� ����������U��EV�u+����� ~P�EVP�����^]� SW�~��$    ��;�t"�;H�}�X��P��X��X�H��P����;�uރ�;}u�_[^]� ���������U��Q���3ŉE��U;Ut>SVW��$    �2�B���;0}�z�����X�Y����;0|�1�y��;Uu�_^[�M�3��v  ��]� ������������U��QS�]W�}��+ǃ���M�=   ��   V�} t{�M��+����+���4ǍǉE�C�;�};�|;�}	�C��;�}���
;��C�|�E�MPSWQ�M��)����U�M�R���ESVP�u�����+������   �^_[��]� �MSWQ�M��o���^_[��]� ������U��SV�uW�}�ٍ�3ɉU�ƃ�t�I ��A��u��	PRWS�M�	����� ~&��   VWS�M�����MQVS�M�u���_^[]� �E;�tPWS�M�����_^[]� �����h��Ph�f �@/  ���������������U���Vh��h�   h�f ���/  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh��h�   h�f ���.  ����t���   ��t�M�UQ�MRQ����^]� U���Vh��h�   h�f ���C.  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh��h�   h�f ���-  ����t���   ��t�M�UQ�MRQ����^]� U��Qh��h�   h�f �x-  ����t���   �E���t�EP�U�����]���f��]�������������U���h��h�   h�f �&-  3Ƀ�;�tK9��   tC�E���   ���M��$Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]ËE�   � �  �P�P�H�H�H��]��U��h��h�   h�f �,  ����t���   ��t]��]����U��h��h�   h�f �i,  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h��h�   h�f �	,  ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h��h�   h�f �+  ����t���   ��t]��3�]��U���Vh��h�   h�f �u+  ����tZ���   ��tP�M�UWQR�M�Q�Ћ���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]á���H�u�QV�҃���^��]����������h��h�   h�f ��*  ����t���   ��t��3��������U��h��h�   h�f �*  ����t���   ��t]��]����U��VWh��h�   h�f �w*  ������tb���    tY�E �M�UP���Q�HR�Q����V�ҡ���H�A�UVR�Ћ��   ���ы�����B�P�MQ�҃� ��_^]á���H�A�UR�Ѓ�_3�^]���U��VWh��h�   h�f ��)  ������tb���    tY�E �M�UP���Q�HR�Q����V�ҡ���H�A�UVR�Ћ��   ���ы�����B�P�MQ�҃� ��_^]á���H�A�UR�Ѓ�_3�^]���U���Vh��h�   h�f �5)  ����tZ���   ��tP�M�UWQR�M�Q�Ћ���u���B�HV�ы���B�HVW�ы���B�P�M�Q�҃�_��^��]á���H�u�QV�҃���^��]����������U���Vh��h�   h�f �(  ����tS���   ��tI�MWQ�U�R�Ћu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]Ë���Q�u�BV�Ѓ���^��]����������������U���Vh��h�   h�f ��'  ����tS���   ��tI�MWQ�U�R�Ћu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]Ë���Q�u�BV�Ѓ���^��]����������������U��h��h�   h�f �Y'  ����t���   ��t]��]����U��h��h�   h�f �)'  ����t���   ��t]��]����U��M��U+u&�A+Bu�A+Bu�A+Bu�A+Bu�A+B]����������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���h���   h�   h�f �E��  �E��E��E�    �E�    �E�    �$  ����t���   ��t	�M�Q�Ѓ�h��h�   h�f �$  ����t���   ��t�UR�M�Q�Ѓ���]ËE�U�M��U��H�M�P�U��H�M��P�H��]������U��E��u����MP�EPQ�C�����]��������������̋�3ɉ�H�H�H�U��V��~ W�}u0jh0pj;j��������t
W���A����3��F��u_^]� �~ t3�9_��^]� ����H<�W�҃�3Ʌ����_�F   ^��]� �����V���F   ����H<�Q��3Ʌ����^��������������̃y t�   ËA��uË���R<P��JP�у��������U����u����H�]� ����J<�URP�A�Ѓ�]� ���������������U������u����H�]Ë���J<�URP�A�Ѓ�]�U������$V��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�SP�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���[t.����B�u�HV�ы���B�P�M�Q�҃���^��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^��]���������������U������$SV��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���t/����B�u�HV�ы���B�P�M�Q�҃���^[��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у����3�������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^[��]����������������U������$SV��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���t/����B�u�HV�ы���B�P�M�Q�҃���^[��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у����3�������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у������������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^[��]��U������$SV��u����H�1�����J<�URP�A�Ѓ�������Q�J�E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@�� j �M�Q�U�R�M��Ћ���Q�J���E�P���у���t/����B�u�HV�ы���B�P�M�Q�҃���^[��]á���P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у����3�������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у������������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�A�U�R�Ћ���Q�Jj j��E�htpP�ы���B�@@��j �M�Q�U�R�M��Ћ���Q�J���E�P���у������������P�E��RHjP�M��ҡ���P�E�M��RLj�j�PQ�M��ҡ���H�u�QV�ҡ���H�A�U�VR�Ћ���Q�J�E�P�у���^[��]����U�졸��H<�A]����������������̡���H<�Q�����V��~ u>���t����Q<P�B�Ѓ��    W�~��t������W�T������F    _^��������U���V�E�P���n�����P�������M���Y�����^��]��̃=�� uK�����t����Q<P�B�Ѓ����    �����tV������V����������    ^������������U���H����H�AS�U�V3�R�]��Ћ���Q�JSj��E�hxpP�ы���B<�P�M�Q�ҋ���H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��  �M�Q�U�R�M��X  ���&  W�}�}���   ������   �U��ATR�Ћ�������   ����Q�J�E�P���ы���B���   ���M�Qj�U�R���Ћ���Q�J���E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Bx��W�M����E���t�E� ��t����Q�J�E�P����у���t����B�P�M�Q����҃��}� u"�E�P�M�Q�M��C  ��������E�_^[��]ËU��U�_�E�^[��]��U���DSV�u3ۉ]�;�u_����H�A�U�R�Ћ���Q�JSj��E�hxpP�ы���B<�P�M�Q�ҋ���H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��A  �M�Q�U�R�M��  ���p  W�}��I �E����   ������   �U��ATR�Ћ�������   ����Q�J�E�P���ы���B���   ���M�Qj�U�R���Ћ���Q�J���E�P�ы���B�P�M�QV�ҡ���H�A�U�R�Ћ���Q�Bx��W�M����E��t�E ��t����Q�J�E�P����у���t����B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*������   P�BH�Ћ���Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��2  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��  �EP�M�Q�M�u��u��  ����   �u���E���tA��t<��uZ������   �M�PHQ�ҋ���Q���ȋBxV�Ѕ�u-�   ^��]Ë�����   �E�JTP��VP�[�������uӍUR�E�P�M��T  ��u�3�^��]����������V��~ u>���t����Q<P�B�Ѓ��    W�~��t������W�Ծ�����F    _^�������̋�� �p����������p���������̅�t��j�����̡���P��  �ࡸ��P��(  ��U�졸��P��   ��V�E�P�ҋuP���J����M�肿����^��]� ��������̡���P��$  ��U�졸��H��  ]��������������U�졸��H���  ]�������������̡���H��  ��U�졸��H���  ]��������������U�졸��H��x  ]��������������U�졸��H��|  ]�������������̡���H��d  ��U�졸��H��p  ]��������������U�졸��H��t  ]��������������U���EV����pt	V��������^]� �������������̸   � �������̸   @� �������̸   � �������̸   � ��������U�졸��H�QV�uV�҃���^]� �3�� �����������3�� �����������3�� �����������U����   h�   ��@���j P��V  �M�Eh�   ��@���R�M��MPQjǅ`���    ��q���� ��]���U����   V�u��u3�^��]�h�   ��@���j P�V  �M�U�Eh�   �M���@���Q�U��U��@����ERPj��`���ǅD�����E�P��E�0��E�p��E�@��E�`��E� ��E�`��E�P��=q���� ^��]������U���   SV�u(3ۉ]���u����H�A�UR�Ѓ�^3�[��]Ë���Q�B<W�M3��Ѕ��N  ��1  �E�����   �MQ�M�赻������B�P�M�Q�ҡ���H�AWj��U�h�pR�Ѓ��M�Q�M��{����u�Wj��U�R�E�P��\���Q�_?�������P��x���R�ο����P�E�P�������P����2  �E���t�E� �� t�M����虻����t��x������膻����t��\�������s�����t�M̃���c�����t����Q�J�E�P����у���t�M��9����}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R�0  ����E$�M�UVP�Ej QRP������������Q�J�EP�у���_^[��]��������̋�`����������̋�` ����������̋�`����������̋�`����������̋�`����������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V����.  �����   �ESP�M��ȸ������Q�J�E�P�ы���B�Pj j��M�h�pQ�҃��E�P�M�茸��j j��M�Q�U�R��d���P�������P�M�Q������P�U�R�ڼ�����P�0  ���M���������M�蹸����d���许���M�覸������H�A�U�R�Ѓ��M�芸����[t	V�.  ����^��]� ���U��EVP����8  �����^]� �����Q��-  Y���������U��E�M�U�H4�M�P �U��M�@��@8P��@<`��@@P��@D0��@Hp��@L ��@P@��@l��@Xp��@\��@`@��@d ��@T`��@h0��@pШ�@t��P0�H(�@,    ]��������������U���   h�   ��`���j P��P  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj��k����8��]��������������̋�`<����������̋�`0����������̋�`@����������̋�`����������̋�`$����������̋�`4����������̋�`(����������̋�`8����������̋�`����������̋�`����������̋�`,�����������U��EHu�E�M�������   ]� �������������U��EHV����   �$����   ^]á��@�����uQ�EP������=�6  }�����^]Ëu��t�jh�pjmj��������t �����������tV��菹���   ^]����    �   ^]ËM�UQR������������H^]�^]飠�����u.�Ơ���!��������t���`���V���������    �   ^]Ã��^]ÍI Щf�m�ȩ��K�����U���EV���V��������Au����H��0  h0qj,�����^��^]� �����U���W������G���U���o������A�  ������A��   ��q������AuR������AuKV����n  ����n  �ȅ�u��^����__��]Ëƙ����ʅ�u�u��E�^������__��]���������Au������=xq��������Au6�����������U������G�����_��������Au�����U����_�
����������Mp  �E����U���l��������A{���������__��]�������������__��]����U����qV�E��������At����q������Au�������m����l�$�l  �����m���^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3�����l;���W���$���!l  ��E����l�$�l  �V����������Au����H��0  h0qj�����^����_u������������^]� ���U������EV�ы�������z!����؋H��0  h0qj5�����U������$�yk  �]��F�$�kk  �}��$�`k  ��E�$�Sk  �^�����&���^��]� ���������������U�졸����   �BXQ�Ѓ���u]� ����Q|�M�RQ�MQP�҃�]� ���U�졸����   �BXQ�Ѓ���u]� ����Q|�M�R8Q�MQP�҃�]� ���U��EV��j �����Qj j P�B�ЉF����^]� ��̡��Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ����Q�MP�EP�Q�JP�у��F�   ^]� ����U��M��P]����U��M��P]����U��M��P]����V����q�F    ����HP�h@�Vh0�h ��҉F����^����������̃y ��qu����PP�A�JP��Y��U��A��u]� ����QP�M�Rj Q�MQP�҃�]� ��U��A��t����QP�M�RQP�҃�]� ������������U��A��t����QP�M�RQP�҃�]� �����������̡���HP���   ��U�졸��HP���   ]�������������̡���HP�QP�����U�졸��HP�AT]����������������̋��     �@    �V����t)����QPP�BL�Ћ���QP��J<P�у��    ^�������������U��SV�ً3�W;�t����QPP�B<�Ѓ��3�s�}�Eh@�W�C����QP�J8h0�h �P�EP�у��9u~M�I ���z u!���@   ����QP���H�RQ�҃�����HP��A@VR�Ћ�F���A;u|�3�9_^��[]� ��������U��SVW��3�9w~<�]����HP��A@VR�Ѓ���t-����QPj SjP�B�Ѓ���tF;w|�_^�   []� ����QP��JLP�у�_^3�[]� �����������̡���PP��JDP�у�������������̡���PP��JHP��Y��������������̡���PP��JLP��Y���������������U��U�E�@R�URP�I���]� �����U��V��~ ��qu����HP�V�AR�Ѓ��Et	V�Ϋ������^]� ����U��E�M�UP��P�EjP�Cf����]��������������̸   �����������U��V�u��t���u6�EjP�Df������u3�^]Ë��1g����t���t��U3�;P��I#�^]������������P�P�P�P �P(�P0�P8�P@�PH�PP�PX����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH������������Dz�u�؋��3�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�����U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A�A �A�A(��l����������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E������X�X]� ̋�3ɉ�H�H�H�V��V藥���FP莥��3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}��+	  S�]����  ��؋���M�U��>���U�@�U���� �U��@�@�B�@�������@���@�   ���]��E��U�;���  �w�����  �w�������F�ݍB��   �U����������������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]����]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]��]��U���E��U��R�э����N�B���B�P���R���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]�����B���B���U����E��������]��E����E����������E������E��E��U����E��]����E��U��E��U��P����E�̋U���������������;���   �ލ���+�������̋�@�������O�]��@���]��@���U������M������]��E��E����E������E����������E��E��U����E��]����E��U��E��E��U�u�����������������������[�[�E���������������a  ��������������Dz���������E��-������������������M����M��E��������������������[H���[P�[X�E����E���������zu������������zh�����CP���CX���CH���CX�������cH���[���[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@��   ������������z]�CX���CP�����cH�CH���CP�������[�[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@�]�CP���CX�����CH���CX�����cP���[0���[8�[@�C8�KX�C@�KP���CH�K@�C0�KX���C0�KP�C8�KH�����[�[ �[(��$���SQ�����E��U�   �����}��M������3�3��u��u���|)�A�����B�4�u�0u��u�p��J�u�u�U�E;�}�Q���E���u��U��1���@���K�I�E    ��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���CX�H�D��@�����U���]�� �K��C0�H���@�KH��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���U����n  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������]��E�E����]���E����]��E��M����@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������U��E��]��E��U������������������9M|��[��_��^���؋�]� ���������ʋE�����׋��@�E�Ѝ��K��C0�H���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���CX�H�E@�E���]����E��������������������M����������]��E��E�;��T�����[������_��^��]� �h��Ph_� �P������������������h��jh_� �/�������uË@����U��V�u�> t/h��jh_� ��������t��U�M�@R�Ѓ��    ^]���U��Vh��jh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh��jh_� ����������t�@��t�MQ����^]� 3�^]� �������U��Vh��jh_� ���I�������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��jh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh��j h_� ����������t�@ ��t�MQ����^]� 3�^]� �������U��Vh��j$h_� ���y�������t�@$��t�MQ����^]� 2�^]� �������Vh��j(h_� ���<�������t�@(��t��^��3�^������Vh��j,h_� ����������t�@,��t��^��3�^������U��Vh��j0h_� �����������t�@0��t�MQ����^]� 3�^]� �������U��Vh��j4h_� ����������t�@4��t�M�UQR����^]� ���^]� ��Vh��j8h_� ���\�������t�@8��t��^��3�^������U��Vh��j<h_� ���)�������t�@<��t�MQ����^]� ��������������U��Vh��j@h_� �����������t�@@��t�MQ����^]� ��������������U��Vh��jDh_� ����������t�@D��t�MQ����^]� 3�^]� �������U��Vh��jHh_� ���i�������t�@H��t�MQ����^]� ��������������Vh��jLh_� ���,�������t�@L��t��^��3�^������Vh��jPh_� �����������t�@P��t��^��3�^������Vh��jTh_� �����������t�@T��t��^��^��������Vh��jXh_� ����������t�@X��t��^��^��������Vh��j\h_� ���l�������t�@\��t��^��^��������U��Vh��j`h_� ���9�������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh��jdh_� �����������t�@d��t�M�UQR����^]� 3�^]� ���U��Vh��jhh_� ����������t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh��jlh_� ���i�������t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh��jph_� ����������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh��jth_� �����������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh��jxh_� ����������t�@x��t�M�UQR����^]� 3�^]� ���U��Vh��j|h_� ���Y�������t�@|��t�MQ����^]� 3�^]� �������U��Vh��h�   h_� ����������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h_� �����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh��h�   h_� ���f�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh��h�   h_� ����������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh��h�   h_� ����������t���   ��t�MQ����^]� 3�^]� �U��Vh��h�   h_� ���v�������t���   ��t�MQ����^]� ��������U��Vh��h�   h_� ���6�������t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh��h�   h_� �����������t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E����������M������U�_��^�U�[���U������������������������P  ��������������D�Ez����P�X��]� �������E�����E����X�M��X��]� ��U���@��m�A���E�    �����]��]��]���m�������]��]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P�1����F�@��R�M������~���Q�M������v;�t�v��P�M�������M����M��M�u�_^[�M�UQR�M�������]� �Q3���|�	��t��~�    t@��Ju��3�����������U��QV�u��;�}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��x+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~!V�1�d$ ���   @u	�����t@��Ju�^�����̋QV3���~�	�d$ ����ШtF��Ju��^�����������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%����E���;�}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$�(��E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ���������������U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�����FP�ތ��3����F�F^��U��SV��WV����^S蹌���E3����~�~;�t_����Q���   h�q��jIP�у��;�t9�}��t;����B���   h�q��    jNQ�҃����uV�K�����_^3�[]� �E�~_�F^�   []� ����������U��SV��WV�����^S�	����}3Ƀ��N�N;���   9��   �G;���   ����Q���  h�q��jlP�у����t=� t@�G��t9����Jh�q��    ���  jqR�Ѓ����u�������_^3�[]� �O�N�G���    �F�RPQ��-  �����t�V�O��RQP�-  ��_^�   []� �����������U��SV��WV�����~W�	���3Ƀ��N�N9M��   �E;���   ��    ����H���  h�qh�   S�҃����t=�} tH�E��tA����Q���  h�q��h�   P�у����u�������_^3�[]� �U�V�,�F   ����H���  h�qh�   j�҃����t��M��ESQR�F�,  �E����t �N���QPR�,  ��_^�   []� ��M�_^�   []� �����U��Q�A�E� ��~JS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U���Ou�_^[�E��Ћ�]� �����������U��S�]V��3�W�~���F�F�CV;C��   �T���W�N���3��F�F����Q���   h�qjIj�Ѓ������   ����Q���   h�qjNj�Ѓ����uV�������_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� 谈��W誈��3��F�F����B���   h�qjIj�у����t[����B���   h�qjNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP��������^]� ���������̡���H���   ��U�졸��H���   V�u�R�Ѓ��    ^]����������̡���P���   Q�Ѓ�������������U�졸��P�EPQ���   �у�]� ̡���H�������U�졸��H�AV�u�R�Ѓ��    ^]��������������U�졸��H�AV�u�R�Ѓ��    ^]��������������U�졸��P��Vh�  Q���   �E�P�ы�����   �Q8P�ҋ�����   ��U�R�Ѓ���^��]��������������̡���P�BQ�Ѓ����������������U�졸��P�EPQ�J\�у�]� ����U�졸��P�EP�EP�EP�EP�EPQ���   �у�]� �U�졸��P�EP�EP�EP�EPQ�JX�у�]� �������̡���P�B Q��Y�U�졸��P�EP�EP�EP�EPQ���   �у�]� �����U�졸��P�EP�EP�EPQ�J�у�]� ������������U�졸��H��   ]��������������U�졸��P�R$]�����������������U�졸��P��x  ]�������������̡���P��|  ��U�졸��P�EP�EP�EP�EPQ�J(�у�]� ��������U�졸��P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U�졸��P�EP�EP�EP�EPQ�J,�у�]� ��������U�졸�V��H�QWV�ҍx�����H�QV�ҋ���Q�M�R4Q�MQ�MQWHPj j V�҃�(_^]� ���������������U�졸��P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U�졸��P�EP�EPQ�J@�у�]� U�졸��P�EPQ�JD�у�]� ���̡���P�BLQ�Ѓ���������������̡���P�BLQ�Ѓ���������������̡���P�BPQ�Ѓ����������������U�졸��P�EPQ�JT�у�]� ����U�졸��P�EPQ�JT�у�]� ����U�졸��P�EP�EPQ���   �у�]� �������������U�졸��P�E���   ��VP�EPQ�M�Q�ҋu�    �F    ������   j P�BV�Ћ�����   �
�E�P�у� ��^��]� ������̡���P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡���H�������U�졸��H�AV�u�R�Ѓ��    ^]��������������U�졸��P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U�졸��P�EPQ�J�у�]� ���̡���P�BQ��Y�U�졸��P�EP�EPQ�J�у�]� U��VW���4����M�U�x@�EPQR�������H ���_^]� �U��VW�������M�U�xD�EPQR��������H ���_^]� �V��������xH u3�^�W��������΍xH�����H �_^�����U��V�������xL u3�^]� W�������M�U�xL�EPQR���z����H ���_^]� �������������U��V���U����xP u���^]� W���?����M�U�xP�EP�EQRP���%����H ���_^]� ��������U��V�������xT u���^]� W��������M�xT�EPQ��������H ���_^]� U��V��������xX u���^]� W�������xX�EP�������H ���_^]� ����U���S�]VW���t.�M���������o����xL�E�P���a����H ��ҍM��0����}��tZ����H�A�U�R�Ћ���Q�J�E�WP�ы���B�P�M�Q�҃����	����@@��t����QWP�B�Ѓ�_^[��]� ������U��V��������x` u
� }  ^]� W�������x`�EP�������H ���_^]� ��U��VW�������xH�EP�������H ���_^]� ���������U��SVW���c����x` u� }  �#���O����x`�E���P���<����H ��ҋ�����H�]�QS�҃�;�A����H�QS�҃�;�,��������M�U�xD�EPQSR��������H ���_^[]� _^�����[]� ��������������U��V�������xP u
�����^]� W�������M�U�xP�EP�EQ�MR�UPQR���{����H ���_^]� ��������������U��V���U����xT u
�����^]� W���=����M�xT�EPQ���+����H ���_^]� ��������������U��V�������xX tW��������xX�EP�������H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u���	  ����t.�E�;�t'����J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡���H��   ��U�졸��H��$  V�u�R�Ѓ��    ^]�����������U�졸��UV��H��(  VR�Ѓ���^]� �����������U�졸��P�EQ��,  P�у�]� �U�졸��P�EQ��,  P�у����@]� �����������̡���H��0  �⡸��H��4  �⡸��H��p  �⡸��H��t  ��U��E��t�@�3�����RP��8  Q�Ѓ�]� �����U�졸��P�EPQ��<  �у�]� �U�졸��P�EP�EP�EPQ��@  �у�]� ���������U�졸��P�EP�EPQ��D  �у�]� �������������U�졸��P�EPQ��H  �у�]� �U�졸��P�E��L  ��VWPQ�M�Q�ҋu������H�QV�ҡ���H�QVW�ҡ���H�A�U�R�Ѓ�_��^��]� ��������������̡���P��T  Q�Ѓ�������������U�졸��P�EPQ��l  �у�]� ̡���P��P  Q�Ѓ�������������U�졸��P�EPQ��X  �у�]� ̡���H��\  ��U�졸��H��`  V�u�R�Ѓ��    ^]�����������U�졸��P�EP�EP�EP�EP�EPQ��d  �у�]� �U�졸��P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���O��z����3��G �G$�G(�G,�G0�G4�G8�G<�G@�GD�GH�GL�GP�GT�GX�G\�_p��G`�Gd�Gh�Gx�����G|   ��_^����������������V��W�>��t7�������xP t$S���q���j j �XPj�FP���]����H ���[�    �~` t����H�V`�AR�Ѓ��F`    _^������������U��SV��Fx����Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR��3������u#���h�r����H��0  h  �҃��E�~P���,~���j j jW�����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ����Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��QV��~d tg�E;Fxt_�N`W�>�M����˹���xP u����(S��踹���UR�XP�E�Pj�NQ��蠹���H ���[�F|_��u�E�Fx�E��t�    �F`^��]� �M�Fx������t�3�^��]� ���������jh�rh�   h�   �w������t���,���3�����������V�������N^��x�����������������U��QS�]VW3��{�����H�QhV�҃������u#�H��0  h�rh�  �҃�_^3�[��]� �}�H�U�R�U�EP���   RV�Ѓ���t�9}�~#�M�<� �4�tj���F  ��t��G;}�|ݍEP��t����_^�   [��]� ��������������U��QS�]VW3��{�����H�QhV�҃������u#�H��0  h�rh�  �҃�_^3�[��]� �}�H�U�R�U�EP���   RV�Ѓ���tӋE;�t�3�9}�~?��E�<� t.������QP�Bh�Ѓ���t�M�<�j���_   ��t�8F;u�|ÍUR�t����_^�   [��]� ���������U��VW�}�7��t�������N�w��V��u�����    _^]�U��USV��F�����N;�~w��@�+�W������%  �yH���@u��u	�   +������J�h(rh�   ��    RP��  �ЋN����t�~_��^^��[]� _�N^[]� �^^[]� ����h��Ph�f �������������������U��h��jh�f �l�������t
�@��t]�����]�������U��Vh��jh�f �;���������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�u���E�NP�у�4�M���u����^]ÍM�u�����^]��U��h��jh�f ���������t
�@��t]��3�]��������U��h��jh�f ��������t
�@��t]��3�]Ë�U���V�u��u�!;  �@�E���:  ���E�F�}� �E�u�E�H�����   �� ��   S�]W�   ;�s��uS��4  Y��u�   �F�Xt}��u�]��}��94  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPW�u�j �3  ��$��u������E�t	�M����_[^�Ë�U��V�:  �@�u���9  jh   �F�m:  YY�F��th   �w3  P�v�7  ���F   ��]3  �f �F��^]Ë�Wh�����`��uV���V�z  ��Y��X�|�^��_�h��� `��yV���V�^  ��Y��X�|�^Ë�U��EV����}k���P�@  Y��^]� ���}k���P�3  YËI�Y�����t�j���Ë�U��j�0#��Y��t�\���M�H�3��\�]Ë�U��E���t������t�j���]Ë�U��Qj �M��Q���h`�������%`� Y�M��_����á`�Ë�U��=�� uh�����  Y�E�`�]�j�cR�9  j �M�������}�e� �w��GN���8 t��p�����t�j�����u��w�  �M��Y�M��������9  �j�cR�_9  j �M������e� ���� �Σ\�����V�#"��Y�\���u��M���M������9  Ë�U��E�@��t
Pj �PD  YY]Ë�U��V��W�};�t>��tP��  Y�& ��t,�? ��t@�8 u�+�S�XS�(*  Y���tSWP�  ��[_��^]� ��U��j j ��C  YY��u�cV�uP�N�����} t�uj �C  YY��u��rP�N�^���^]Ë�U��V��M3��N�N�F   ��r�F�F�Fh�r��A�#�����^]� j��R�8  ��u���rV�E�   �/����FY��tP�  Y�f ��f�E8  Ë�U��V�������EtV� ��Y��^]� j�cR�7  �`�3���;�unV�M�������`��u���;�uKj �M ��Y;�t
V��������V���w����N�F?   �$�r�T����Ή5d������d��|��M���M��������7  Ë�U��Q�E;Pu�	;u3�@�3�]� ��U��E�U��H]� ��U��QQ�u��u�U�R�P�������� ��U��E;Hu� ;Eu3�@�3�]� �AËAø��Ë�U���EV����rtV�x��Y��^]� ��U��Q�u�e� ��C  Y�MP��E���E�� ��U��Q�e� �}uhds�
�u��C  YP�M�E���E�� ��U��VW���w,��vW�u�V�6����u�_^]� ��VWj ��������F(��t�8P����Y�ǅ�u�F,�f( ��t�8P����Y�ǅ�u�f, _^Ë�U��V�u�~ v�F������8 �������v0��t��辱��V�x��Y^]���  ��U��V�u���  ��s��^]� ��U����E�E�EP�M��D  hи�E�P�E��s�  ̋�U��V�u����  ��s��^]� ��U����E�E�EP�M���  h��E�P�E��s�=  ̋�U��V�u���}  ��s��^]� ��U��V���  �EtV���Y��^]� ��U���V�u��u�A3  �@�E��3  ���E�F�}� �E�u�E�H�����   �� ��   S�]��   s!��uS�w-  Y��u�   �F�X��   ��u�]��}��W,  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPh   �u�j �+  ��$��u������E�t	�M����[^�Ë�Vj���Y��P��  YY��^Ë�V���6��   �6�X��YY^��1��   Y��1�  YË�U���u�E�4��s�u�%A  ��]Ë�U��MS3��ًу���   @V��@t���t����;���3�;�t��tF��u��<�t u3��U��t"��
t�uj �u�|�������t	P�y  Y���uV�u�`���������t���tjj V��A  ����tV�ˋ�^[]Ë�U��]�M�����U���u�(`]Ë�U���u�,`]Ë�U���u�0`]Ë�U���u�4`]Ë�U��= � u]��A  �u� ��8`� �����]��� ������ �P�<`��t�Ѓ= �
r����̋L$WSV��|$��to�q��tU���L$���:�t��t���:�t
��u�^[_3�Ê��:�u�~��a��t(���:�u��A��t�f���:�t��3�^[_���A  �G�^[_Ë�^[_Ë�Q�Xt�*B  YË�U��V��������EtV�!��Y��^]� ��U��E��	Q��	P�dB  ��Y�Y@]� ��U��E��t���8��  uP�	  Y]Ë�U��EV���F ��uc�vN  �F�Hl��Hh�N�;��t����Hpu�%L  ��F;��t�F����Hpu�D  �F�F�@pu�Hp�F�
���@�F��^]� ��U������3ŉE�V��u�S  j^�0�R  �7  �uW�Q  YY;Er� �׋�H��u"�? ��t�<a|<z, �A�9 u�3���   j�p�   j j j�WVQS��'  �ȃ�$�M��u�R  � *   �R  � �   9Ms� �~R  j"�c�����~Ej�3�X���r9�A=   w�R  �ą�t� ��  �P��   Y��t	� ��  ���M�E���e� �}� u�R  �    뀋j�pQ�u�j�WV�pS� '  ��$��t�u��uW��   �������Q  j*Y����u������Y�ƍe�^�M�3��
  �Ë�U���SW�u�M�������u�}�]��i����}� Y_[t�M��ap��Ë�U��j �u�u������]Ë�U��=,� u;�E��u�XQ  �    ��P  3�]À8 ��t+�
��a|
��z�� �
B�: u�]�j j��u�_����E��]Ë�U��UVW��t�}��u��P  j^�0�P  ���3�E��u����+���@��tOu��u� ��P  j"Y�����3�_^]�;��u���#Q  ������̋T$�L$��ti3��D$��u���   r�= � t��Q  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$ø�V�`��d��M�h��M�l��M�p�BM�t��x�nV�|�^M����L���LLË�U�������} t��\  ��]��������������U��WV�u�M�}�����;�v;���  ���   r�= � tWV����;�^_u��\  ��   u������r)��$����Ǻ   ��r����$����$�����$�d���� �D�#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I �����������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�l������$���I �Ǻ   ��r��+��$�p��$�l���������F#шG��������r�����$�l��I �F#шG�F���G������r�����$�l���F#шG�F�G�F���G�������V�������$�l��I  �(�0�8�@�H�P�c��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�l���|��������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�ËA��u�ltË�U��} W��t-V�u�6  �pV�  YY�G��t�uVP��������G^_]� ��V��~ t	�v�,  Y�f �F ^Ë�U��EV��f �dt�F �0������^]� ��U��V�uW��;�t�����~ t�v���V�����F�G��_^]� �dt�{�����U��V�EP��������t��^]� ��U��V���dt�J����EtV�P��Y��^]� ��U��V�u��f �dt�F �]�����^]� ��U��V�u���������t��^]� ����������������������U��WV�u�M�}�����;�v;���  ���   r�= � tWV����;�^_u��W  ��   u������r)��$�� �Ǻ   ��r����$����$�� ��$�4 ����� #ъ��F�G�F���G������r���$�� �I #ъ��F���G������r���$�� �#ъ���������r���$�� �I � � | t l d \ T �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�� ��� � � � �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�<�����$���I �Ǻ   ��r��+��$�@�$�<�Pt��F#шG��������r�����$�<�I �F#шG�F���G������r�����$�<��F#шG�F�G�F���G�������V�������$�<�I ��  3�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�<��LTdx�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_����������������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[Ë�U��} t-�uj �5���D`��uV�F  ���@`P�=F  Y�^]Ë�U��� �EVWjY��t�}��E��E_�E�^��t� t�E� @��E�P�u��u��u��H`�� jhH��X  3��}�3��u;���;�u�	F  �    �E  ����   V��  Y�}��F@uoV�3X  Y���t���t�����ȃ���� ������A$u)���t���t��������� ������@$�t�E  �    �)E  �M��9}�u�Nx
��A��V��S  Y�E��E������   �E��
X  ËuV�  Y�jhh��W  3��}�3��u;���;�u�E  �    �D  ����   V��  Y�}��F@uoV�?W  Y���t���t�����ȃ���� ������A$u)���t���t��������� ������@$�t�D  �    �5D  �M��9}�u!�Nx��E�����V�u��X  YY�E��E������   �E��W  ËuV�  YË�U��SV�uW����F@uoV�vV  Y���;�t���t�ȃ�������� �����A$u%;�t���t�ȃ������ �����@$�t��C  �    �oC  ��_^[]Ë];�t�F�u��y�u�~ uV�kY  Y�;Fu	�~ u�@���F@�t	8t@�볈�F�F�����F��%�   �jh����U  3�9E����u�=C  �    ��B  ����,�u�  Y�e� �u�u�����YY�E��E������	   �E���U  ��u�L  Yø��á@
Vj^��u�   �;�}�ƣ@
jP�  YY�(���ujV�5@
��  YY�(���ujX^�3ҹ����(���� ����@�|�j�^3ҹ��W������ �����������t;�t��u�1�� B��0�|�_3�^���  �=�� t�CX  �5(��i���YË�U��V�u���;�r"�� �w��+�����Q��\  �N �  Y�
�� V�0`^]Ë�U��E��}��P�\  �E�H �  Y]ËE�� P�0`]Ë�U��E���;�r= �w�`���+�����P�[  Y]Ã� P�4`]Ë�U��M�E��}�`�����Q�j[  Y]Ã� P�4`]Ë�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�[S  YP�)c  ��;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV��R  P�c  Y��Y��3�^]�jh��� S  3��}�}�j�i[  Y�}�3��u�;5@
��   �(���98t^� �@�tVPV�h���YY3�B�U��(����H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u�(��4�V�q���YY��E������   �}�E�t�E��R  �j��Y  Y�jhй�&R  3�9uu	V����Y�'�u�t���Y�u��u����Y�E��E������	   �E��/R  ��u����Y�j�����Y�jh���Q  �e� 3��u������u�3?  �    ��>  ����   �]��t	��t��@uׅ�t��@u�}�G�=���v뿋}����uV�����Y�e� V����V�b  YY�f�����N��t���Fj_�-�E��u W�  Y��u���M����N  �	��   �N�~�F��f �E������	   �E��0Q  ��u����YË�U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$����U��QQSVWd�5    �u��E�j �u�u��u�PD �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�m  �� �E�_^[�E���]Ë�U��V��u�N3������j V�v�vj �u�v�u�hm  �� ^]Ë�U���8S�}#  u�A�M�3�@�   �e� �E�m����M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E��7  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M������E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u�2l  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����+���u��l  �MN��k�E�9H};H~���u	�M�]�u�} }̋EF�0�E�;_w;�v�l  ��k�E�_^[�Ë�U��EV�u��C6  ���   �F�56  ���   ��^]Ë�U��� 6  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V��5  �u;��   u��5  �N���   ^]���5  ���   �	�H;�t���x u�^]�l  �N�H�ҋ�U�������e� �M�3��M�E��E�E�E@�E�c�M��E�d�    �E�E�d�    �uQ�u�l  �ȋE�d�    ���Ë�U��V�u��u3��a�} u�`:  j^�0�:  ���H�} t9urV�u�u�k��������uj �u�������} t�9us�:  j"Y����jX^]Ë�U���SVW�}��t�} t�u��u��9  �    �9  3�_^[�ËM��t���3���9Ew��}�F  �M��}��t�F�E���E�   ����   �N��  t/�F��t(��   ��;�r��W�u��6����)~>��+�}��O;]�rO��tV����Y��u}�}� ��t	3ҋ��u�+�W�u�V�|K  YP�J[  �����ta��;�w��M�+�;�rP�}��)�E�� VP�fM  YY���t)�E��FK�E����E�   ���A����E������N ��+�3��u������N �E���jh��$K  3�9ut!9ut3�9u��;�u�8  �    �*8  3��:K  ��u�R���Y�u��u�u�u�u�P������E��E������   �E����u����YË�U��} u�&8  �    ��7  ���]�V�u��u�	8  �    �7  �����u�m  Y�ȉ#ʃ���V;�t3�^]Ë�U��V�u�FW��ty�}��t
��t��uh���F��uV�ti  EYU3�V�]����FY��y����F��t�t�   u�F   W�u�uV�I  YP�gm  #����t3���L7  �    ���_^]�jh0��I  3�9E����u�"7  �    ��6  ����B�u��t
��t��u��u�����Y�e� V�u�u�u�
������E��E������	   �E��I  ��u����YË�U��} u�6  �    �S6  ���]ËE��t�j �p�0�u�K�����]Ë�U��V�uW�����u�o6  �    �6  ��D�F�t8V����V���!Z  V�H  P��m  ����y�����F��tP�t����f Y�f ��_^]�jhP��H  �M��3��u������u��5  �    �5  �����F@t�f �E��H  �V����Y�e� V�<���Y�E��E������   �ԋuV�����YË�U���u�P`��u�@`�3���tP�5  Y���]�3�]Ë�U��� �e� WjY3��}��_��u�S5  �    ��4  �����9Et�V�8  Y�����E�I   �u�u��M�;�w�E��u�E��u�uP�U���Ë�U��V�u�EPj �uh	��v�����^]Ë�U��Q�e� S�]��u3��   V��ru�s���tn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9u�r��.�@��I��F�@��I��<�@��I��2�@��I��(�M�E�u�����t:u@FA;�r�3�^[��� �	+����U��j
j �u�K  ��]��5H��<`��t��j�~  jj ��   ����   jhp��XF  �E��uz�2B  ��u3��8  �G0  ��u�7B  ��蟆  �X`�$����  ���LC  ��y��,  ���#�  ��x 褂  ��xj ��J  Y��u����   �XE  ��3�;�u[9=�~����}�9=��u�L  9}u�(E  �,  �A  �E������   �   3�9}u�=���t�c,  ��j��uY�",  h  j�)  YY��;�����V�5���5\��<`�Ѕ�tWV�[,  YY�T`��N��V�����Y�������uW�.  Y3�@�HE  � jh����D  ����]3�@�E��u9���   �e� ;�t��u.��t��tWVS�ЉE�}� ��   WVS�C����E����   WVS蔑���E��u$��u WPS耑��Wj S������t��tWj S�Ѕ�t��u&WVS�������u!E�}� t��t��tWVS�ЉE��E������E���E��	PQ�)�  YYËe��E�����3��PD  Ë�U��}u�$�  �u�M�U�����Y]� ��U��S�]���woVW�=�� u�~  j��|  h�   �H  YY��t���3�@Pj �5���\`����u&j^9\�tS�Y�  Y��u����0  �0��0  �0��_^�S�8�  Y��0  �    3�[]���̃=�� ��  ���\$�D$%�  =�  u�<$f�$f��f���d$��  � �~D$f(�tf(�f(�fs�4f~�fT�tf��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$蒅  ���D$��~D$f��f(�f��=�  |!=2  �fT�t�\�f�L$�D$����f��tfV�tfT�tf�\$�D$���������������̃= � t-U�������$�,$�Ã= � t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$�Ë�U��QSV�5<`W�5 ����5���؉]��֋�;���   ��+��G��ruS讈  �؍GY;�sH�   ;�s���;�rP�u��'  YY��u�C;�r>P�u��  YY��t/��P�4��8`� ��u�=8`�׉��V�ף���E�3�_^[�Ë�Vjj �}
  YY��V�8`� ������ujX^Ã& 3�^�jh���@  ��D  �e� �u�����Y�E��E������	   �E��@  ���D  Ë�U���u���������YH]�����������̺ u�Q�  � u�̇  ���������z�����������������̃��$�݌  �   ��ÍT$舌  R��<$�D$tQf�<$t�@�  �   �u���=� ���  �   �@�鰌  �  �u,��� u%�|$ u����  �"��� u�|$ u�%   �t����-0��   �=� �V�  �   �@��_�  ZË�U������3ŉE��US3�VW;�~�E��I8t@;�u������+�H;�}@�E�]�9]$u�E� �@�E$�5h`3�9](SS�u���u��   P�u$�֋��}�;�u3��R  ~Cj�3�X����r7�D?=   w�u,  ��;�t� ��  �P����Y;�t	� ��  ���E���]�9]�t�W�u��u�uj�u$�օ���   �5d`SSW�u��u�u�։E�;���   �   �Mt)�E ;���   9E���   P�uW�u��u�u���   �}�;�~Bj�3�X����r6�D?;�w�+  ��;�th���  ���P�����Y;�t	� ��  �����3�;�t?�u�W�u��u��u�u�օ�t"SS9] uSS��u �u�u�WS�u$�``�E�W�%���Y�u������E�Y�e�_^[�M�3��+����Ë�U����u�M������u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap����i%  �ȋAl;��t����Qpu�##  ���   Ë�U����u�M������E����   ~�E�Pj�u诊  ������   �M�H���}� t�M��ap��Ë�U��=,� u�E����A��]�j �u����YY]Ë�U����u�M��%����E����   ~�E�Pj�u�0�  ������   �M�H���}� t�M��ap��Ë�U��=,� u�E����A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u豉  ������   �M�H���}� t�M��ap��Ë�U��=,� u�E����A��]�j �u����YY]Ë�U����u�M��'����E����   ~�E�Ph�   �u�/�  ������   �M�H%�   �}� t�M��ap��Ë�U��=,� u�E����A%�   ]�j �u�~���YY]Ë�U����u�M������E����   ~�E�Pj�u謈  ������   �M�H���}� t�M��ap��Ë�U��=,� u�E����A��]�j �u����YY]Ë�U���L���3ŉE�S3�V�uW�]ԉ]�]��]؉]܉u��]�9^�  �F9u P�F0h  P�E�SP�u  ������  j�  j��  W�E���  jW�E��  jW�E��  jh  �E��  ��$�E�9]��  9]��v  ;��n  9]��e  9]��\  �Eԉ3��M܈@=   |�E�P�v�l`���2  �}��(  �E�EЃ�~.8]�t)�E�:�t �x�����M�� �G;�~��8X�uڋE�SS�v   Ph   �u܉E�jS蝈  �� ����  �M��E�S�v��   W���   QW@Ph   �vS������$����  �E�S�v�   WP�E�W@Ph   �vS�S�����$���b  �E�}����   3҃}�f��U؉Mč��   �_�Z��M����   �MȈ~U8]�tP�M�M�:�tD�I��҉M�;�(��H   ��M��E� �  f����M̋M��	9M�~�M���M�8Y�u�h�   ��   QP����j��   PW�����E�j��   QP�������   ��$;�tKP� `��u@���   -�   P�������   ��   +�P�w������   +�P�i������   �^������E��    ���   �E����   �Eĉ��   �E����   �Eȉ��   �EЉ��   �u�����Y���o�u��
����u������u�������u������3ۃ�C�ˋ��   ;�tP� `���   ���   ǆ�   Pvǆ�   �zǆ�   X|ǆ�      3��M�_^3�[�������  �ȋAl;��t����Qpu��  �@���  �ȋAl;��t����Qpu�  ��Ë�U��VW3��u������Y��u'9(�vV�$`���  ;(�v��������uʋ�_^]Ë�U��VW3�j �u�u��  ������u'9(�vV�$`���  ;(�v��������uË�_^]Ë�U��VW3��u�u�#�  ��YY��u,9Et'9(�vV�$`���  ;(�v��������u���_^]Ë�U��VW3��u�u�u��  ������u,9Et'9(�vV�$`���  ;(�v��������u���_^]�Pd�5    �D$+d$SVW�(�表�3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(�表�3�P�e��u��E������E�d�    ËM�d�    Y__^[��]QË�V���t��t;�tWj6Y���  P�  Y_^Ë�U��SW3�3�9]~"V�u���6�u�u蘘  ����uG;}|�^_[]�SSSSS�C!  ̋�U��SVW�}h�   3�SW�-����u�����u3���   <.u1�F8t*jP���   jP���  ����u���   ��SSSSS��   h`~V�]臘  ;��   �} �<0�u��@��   ��.t|PVj@�u�;�}u��@sh��_tcP�EVj@��@��}uQ��sL��t��,uCP�EVj��P�d�  ����u4��,�=������5����E�wh`~V���  ��YY�k������_^[]�3�PPPPP�=�����U��SV�uV�u�u������3ۅ�uA�F@8tPhd~j�u�u�g��������   8^[tPh�jj�u�u�E�����]�SSSSS�  ̋�U���S3�ChU  �]��H���Y�E����=  W�x� ��vX�Q  hl~�5�}jSW������FX���E��}�E�hh~SW苖  ������   �E��H�1�M��0�Y  YY��t�e� �E��0�E�hl~�E��E��0jSW�������}��}|��}� uU�FP� `��tP�Ӆ�u	�vP�����Y�FT��tP�Ӆ�u	�vT����Y�E��fT �fL �FP�~H���Z3�PPPPP�  �u������FP�= `3�Y;�tP�ׅ�u	�vP�o���Y�FT;�tP�ׅ�u	�vT�X���Y�Fh�^T�^L�^P�^H_[�Ë�U���   ���3ŉE��ESV�uW�}��d����E��\�����`����  ���   ��T������   ���   K  ��X�����h�������  ��d��� ��  �} ��  �>CuS�~ uMh�r�u��d����A�������u'��tf�f�Gf�G��`�����t�  ��d����C  3�PPPPP�x  V�  ��   Y��P���;�s,V��h����z  YY����   V��X����d  YY����   ��L��� ��l���VP�����YY����   ��l���PSP�F�  ������   �C��T������l���PW��h����������> t
��P���;�r��L����c@PVW��X���讔  �����%���3�9�\���tjS��\����e�����9�`���tj��T�����`����G�������h����u��d������������u��h����VVVVV�����3��M�_^3�[�"����Ë�U����  ���3ŉE��ES��W��p�����h����~  ��S��\���P��P���Ph�   ��x���P��h�����������u3��M�_3�[����������sH��x���P��
  YY��u�CH�Ӎ�x���P�?  ��P��t����5���YY��l�����t��CH��p�����h����D���X���� ��H����Ak��jP��d�����8���P�����F��x���Q��t�����L�����l��������QP���������	  ��l�����X������CH��P����j��P���P��d�����������p����  ��\�����t��� �F���  ���  ��d������  �V;t6���t������d�����@����P�H��@�������t�����d���|��-��t�����t#����  ����  �P���  ���d����H��t���urj�v��x����vPjh�}jj ��|  �� ��t<3���  f!�Ex���@��r�h�   �5P���x���P��  �����@���  ����   �F���  ���  ���   ��p���u	��\����F��p���k�V���}Y��t1��h�����l����CH�l�����H���Y��X������L����F������h�����t.��p�������4�� `��u�4��#����sT�����cL YY��p�����l�������    ���Y���3�PPPPP��  ̋�U���   ���3ŉE��ESV3ۋ�W��h���;�t;�tP����Y��  ɋD�H��  ǅp���   ��t���;���  �8L�0  �xC�&  �x_�  ��hp~W���  ��YY����   +ǉ�p�����   �;;��   ǅl���   ��}���p���PW�6���������u�6��  Y9�p���t��l��������}~�Chh~S诏  ��3�YY;�u	�;;��   ��l���DWS��x���h�   P�Ə  ����uT��l�����h�����=x�����x���P�t���Y��t��t�����? t
G�? ����3�9�t�����   ��h����   VVVVV�g  3��xSSSh�   ��x���QP�������;�t\�~H��t5�7��x���P�V  YY��t��x���P�������Y��u!�p������t���C����~�3�9�p���u9�t���t�3����M�_^3�[�������jhк��)  �e� �}v�e  �    �  3��9  �#  ���u���  �Np�e� 3�GWh�   �x���YY�؉]܅���   j�2  Y�}��Nl�������e� �   �u�M���X���Y�E�����   �} th���u�U  YY��t�=,�j�1  Y�E�   �~lSW�  S�%  ���Fpu?���u6�7h����  YY������   ������   �H����   � ��e� �   �.�]܋u�3�Gj�f0  YËu�j�Z0  Y��S�  S�?  YY�E������   �E���(  Ëu�fp�������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U��V�u��x	胪  ;0|�z�  �0�y�  ��^]Ë�U��SV�  ��3�;�u�x~�"W��   9^$ujW�i���YY�F$;�u
�x~_^[]��u�v$����PWV���������u����SSSSS�@  �jh��W'  3ۉ]�3��};���;�u�  �    �b  3��y3��u;���;�t�3�8��;�t��U�  �E;�u�  �    �ʉ]�8u �r  �    j��E�Ph���\�  ���P�uVW�x�  ���E��E������	   �E���&  ��u����YË�U��V�u�F��u�  �    ����g���}�FuV萯  E�e YV�����FY��y����F��t�t�   u�F   �u�uV�&  YP�u�  3Ƀ�������A�^]�jh(��&  3�9E����u�  �    �#  ����?�u��t
��t��u��u�=���Y�e� V�u�u�������E��E������	   �E���%  ��u�|���Y�蠰  ��tj袰  Y�`�tjh  @j�,  ��j�*,  ̋�U��M�`��U#U��#�ʉ`�]�������������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[�jhH��f$  j��,  Y�e� �u�N��t/�4��0��E��t9u,�H�JP�����Y�v�����Y�f �E������
   �U$  Ë���j�+  Y��̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP����3��ȋ��~�~�~����~����p����F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  ���3ŉE�SW������P�v�l`�   ����   3�������@;�r�����ƅ���� ��t0���������;�w+�@P������j R�O������C����u�j �v�������vPW������Pjj ��q  3�S�v������WPW������PW�vS�������DS�v������WPW������Ph   �vS������$3���E������t�L���������t�L ��������  ���  @;�r��R��  ǅ��������3�)�������������  ЍZ ��w
�L�Q ���w�L �Q����  A;�rƋM�_3�[�!�����jhh��I!  �	  ������Gpt�l t�wh��uj �(  Y���a!  �j�)  Y�e� �wh�u�;5��t6��tV� `��u��p�tV����Y����Gh�5���u�V�`�E������   뎋u�j�R(  YË�U���S3�S�M��d����8����u�8�   �t`8]�tE�M��ap��<���u�8�   �p`�ۃ��u�E��@�8�   ��8]�t�E��`p���[�Ë�U��� ���3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�����   �E��0=�   r����  �t  ����  �h  ��P�x`���V  �E�PW�l`���7  h  �CVP�r���3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�+����M��k�0�u������u��+�F��t)�>����E�����D;�FG;�v�}���> uЋu��E����}��u�r�ǉ{�C   �i���j�C�C����Zf�1f�0����Ju������������L@;�v����~� �0����C��   �@Iu��C�����C�S��s3��ȋ�����{����958��T�������M�_^3�[������jh���@  �M���  ���}�������_h�u�q����E;C�W  h   ����Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh� `��u�Fh=p�tP����Y�^hS�=`���Fp��   �����   j�	&  Y�e� �C�H��C�L��C�P�3��E��}f�LCf�E<�@��3��E�=  }�L����@��3��E�=   }��  ����@���5��� `��u���=p�tP�����Y���S���E������   �0j�$  Y��%���u ��p�tS����Y�G
  �    ��e� �E���  Ã=� uj��V���Y��   3�Ë�U��SV�5`W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{���t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5 `W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{���t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�U��SV�u���   3�W;�to=8�th���   ;�t^9uZ���   ;�t9uP��������   ��z  YY���   ;�t9uP��������   �[x  YY���   ��������   ����YY���   ;�tD9u@���   -�   P�������   ��   +�P�������   +�P�s������   �h��������   =��t9��   uP��s  ���   �?���YY�~P�E   ����t�;�t9uP����Y9_�t�G;�t9uP����Y���Mu�V�����Y_^[]Ë�U��W�}��t;�E��t4V�0;�t(W�8�j���Y��tV������> Yu�� �tV�s���Y��^�3�_]�jh����  �  ����Fpt"�~l t�  �pl��uj �~   Y����  �j�"  Y�e� �5����lV�Y���YY�E��E������   �j��   Y�u��j �8`��|`� ��V�5����`����u�5X��<`��V�5����`��^á�����tP�5`��<`�Ѓ���������tP��`�����    jhȻ��  h���`�u�F\���f 3�G�~�~pƆ�   CƆK  C�Fhp�j�!  Y�e� �vh�`�E������>   j��   Y�}��E�Fl��u����Fl�vl����Y�E������   �  �3�G�uj��  Y�j��  YË�VW�@`�5����������Ћ���uNh  j�������YY��t:V�5���5\��<`�Ѕ�tj V�����YY�T`�N���	V臾��Y3�W��`_��^Ë�V��������uj�v  Y��^�jh��  �u����   �F$��tP�:���Y�F,��tP�,���Y�F4��tP����Y�F<��tP����Y�F@��tP����Y�FD��tP�����Y�FH��tP����Y�F\=��tP�ս��Yj�x  Y�e� �~h��tW� `��u��p�tW訽��Y�E������W   j�?  Y�E�   �~l��t#W����Y;=��t�� �t�? uW�*���Y�E������   V�P���Y��  � �uj�  YËuj�  YË�U��=���tK�} u'V�5���5�`�օ�t�5���5�����ЉE^j �5���5\��<`���u�x���������t	j P��`]Ë�Wh���`����u	�����3�_�V�5�`hD�W��h8�W�T���h,�W�X���h$�W�\��փ=T� �5�`�`�t�=X� t�=\� t��u$��`�X���`�T�.C�5\��`��|`��������   �5X�P�օ���   �  �5T��58`���5X��T����5\��X����5`��\��֣`���  ��tc�=<`h�D�5T����У�����tDh  j������YY��t0V�5���5\����Ѕ�tj V����YY�T`�N��3�@��i���3�^_Ë�U��3�9Ev�M�9 t@A;Er�]Ë�U��E�d�]Ë�U���(  ���3ŉE�S�]W���tS�ܠ  Y������ jL������j P������������������0�����������������������������������������������f������f������f������f������f������f��������������E�M������ǅ0���  �������I��������M�������M��������������`j ����`������P��`��u��u���tS��  Y�M�_3�[�����Ë�Vj� �Vj�������V��`P��`^Ë�U���5d��<`��t]���u�u�u�u�u�����3�PPPPP�������Ë�U��E3�;���tA��-r�H��wjX]Ë���]�D���jY;��#���]��W�����u�X�Ã���D�����u�\�Ã�Ë�U��V������MQ�����Y�������0^]��������Q�L$+ȃ����Y�ڞ  Q�L$+ȃ����Y�Ğ  ��U���(  �p��l��h��d��5`��=\�f���f�|�f�X�f�T�f�%P�f�-L������E �t��E�x��E������������  �x��t��h�	 ��l�   ��������������������`���j��  Yj ��`hP���`�=�� uj�ǝ  Yh	 ���`P��`��f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U���j
��`� �3�Ë�U���V�u�M������u�P�F�  ��e�F�P�d�����Yu��P�)�  Y��xu���M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M��s����E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�d�  �M��E��M��H��EP��  �E�M����Ë�U��j �u�u�u������]Ë�V����tV�7���@PV�V茬����^Ë�U��j �u�d���YY]Ë�U��j �u�����YY]Ë�U���SV�u�M����1���3�;�u"�����j^�0�����}� t�E��`p���^[��9Mv�9M~�E�3���	9Ew	����j"��W8Mt�U3�9M��3Ƀ:-����ˋ��6����}�?-��u�-�s�} ~�N�E�����   � � F�3�8E��E��}�u����+�]hX�SV��������ut�N9Et�E�G�80t/�GHy���F-��d|�jd_�� F��
|�j
_�� F�� F���_t�90uj�APQ�$������}� t�E��`p�3������3�PPPPP�����̋�U���,���3ŉE��ESV�uW�}j[S�M�Q�M�Q�p�0� �  ����u�`�����������m�E��t���u��3Ƀ}�-��+�3Ʌ���+��M�Q�NQP3��}�-��3Ʌ�����Q�<�  ����t� ��u�E�j P�u��V�u��������M�_^3�[�%����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �ۥ��9}}�}�u;�u#����j^�0�$����}� t�E�`p����  9}v؋E��� 9Ew	�J���j"�ȋ}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW�$�������t�}� � ��  �M�ap��  �;-u�-F�} �0����$�x�Fje��V�&�  YY���U  �} ���ɀ����p��@ �;  %   �3��t�-F�]������$�x����0�F�O�����  �3���'3��u$�F0�O����� ���u�U���E��  ��F1����F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~L�W#U���M�#E���� �ٜ  f��0����9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� 膜  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V莦����u�E�8 u���} �4����$�p���W��  3�%�  #�+E�SY�x;�r	�F+����F-������ڋ��0;�|$��  ;�rSQRP��  0�F�U�����;�u��|��drj jdRP�  0��U�F����;�u��|��
rj j
RP蜚  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u���w�ٍM�N�l�����u#����j^�0������}� t�E��`p����   �} v׀} t;uu3��?-���f�0 �?-��u�-�s�G��V�^�����@PVS�����0�������} ~QV�^����@PVS�����E����   � � ������y&�߀} u9}|�}�}������Wj0S跤�����}� t�E��`p�3�_^[�Ë�U���,���3ŉE��EVW�}j^V�M�Q�M�Q�p�0褘  ����u�����0�������lS�]��u������0�������S���;�t3Ƀ}�-����+��u�M�Q�M��QP3��}�-���P�ܖ  ����t� ��u�E�j VS���N�����[�M�_3�^�ˣ���Ë�U���,���3ŉE��EV�uWj_W�M�Q�M�Q�p�0��  ����u�C����8��������   �M��t�S�]�3�K�}�-���<0���u��+ȍE�P�uQW�2�  ����t� �W�E�H;������|-;E}(��t
�G��u��G��u�E�j�u���u��������u�E�jP�u���u�u������[�M�_3�^�ޢ���Ë�U��E��et_��EtZ��fu�u �u�u�u�u�'�����]Ã�at��At�u �u�u�u�u�u������0�u �u�u�u�u�u�o�����u �u�u�u�u�u�o�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3���`��8`��`�����(r�_^Ë�Vh   h   3�V��  ����t
VVVVV�����^�W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����j h   j ��`3Ʌ����������5����`�%�� Ë�U��V�u��u�U����    �������   �F����   �@��   �t�� �F��   ���F�  u	V��  Y��F��v�vV�O  YP�C�  ���F����   �����   �F�uQV�%  Y���t0V�  Y���t$WV�  ��V�<� ���  ��Y��Y_�����@$�<�u�N    �~   u�F�t�   u�F   ��N�A���������	F�f ���^]Ë�U���LV�E�P��`j@j ^V�q���YY3�;�u����  ��   � ��5�;�s6���H��f�@� 
�Hf�@ 
�@!
�H3�H/�5 ���@�P���   ;�r�SWf9M��  �E�;��  ����E�þ   �E�;�|��9�}k�$�j@j �����YY��tQ�� ��   �;�s1���H���` �`��`3 f�@� 
f�@ 

�@/ ���@΍P�;�r҃�9�|����3���~r�E�� ���t\���tW�M��	��tM��uP��`��t=����������4� ��E�� ��E�� �Fh�  �FP��`����   �F�E�G�E�;�|�3ۋ���5 �����t���t�N��q�F���uj�X�
�C�������P��`�����tB��t>W��`��t3%�   �>��u�N@�	��u�Nh�  �FP��`��t,�F�
�N@�����C���h����5���`3�_[^�Ã������VW� ����t6��   ;�s!�p�~� tV�,`���@   �N�;�r��7�����' Y���� �|�_^Ë�U��E��u�����    �?������]Ë@]��������h�\d�5    �D$�l$�l$+�SVW���1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s35��W��E� �E�   �{���t�N�38�1����N�F�38�!����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t��脆  �E���x@G�E��؃��u΀}� t$����t�N�38讛���N�V�3:螛���E�_^[��]��E�    �ɋM�9csm�u)�=�� t h����  ����t�UjR������M�U�$�  �E9Xth��W�Ӌ��&�  �E�M��H����t�N�38�����N�V�3:�����E��H��躅  �����9S�O���h��W���х  ������U��QV�uV������E�FY��u�q���� 	   �N ����/  �@t�V���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�"����� ;�t������@;�u�u蔘  Y��uV��   Y�F  W��   �F�>�H��N+�I�N;�~WP�u��  ���E��M�� �F����y�M���t���t����������� ������@ tjSSQ�z   #����t%�F�M��3�GW�EP�u�v  ���E�9}�t	�N �����E%�   _[^�Ë�U����h   ����Y�M�A��t�I�A   ��I�A�A�A   �A�a �]�jh��X���3ۉ]�j��  Y�]�j_�}�;=@
}T���(�9�tE���@�tP至��Y���t�E��|(�(����� P�,`�(��4�迢��Y�(���G��E������	   �E������j�i  YË�U��hp���`��th`�P��`��t�u��]Ë�U���u�����Y�u��`�j��  Y�j�  YË�V������V�(>  V����V��7  V�Ö  V���  V�'  ��^Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=\t th\t�d�  Y��t
�u�\tY����h�ahta����YY��uTVWh��}����Ha�paY��;�s���t�Ѓ�;�r�=� _^th����  Y��tj jj ��3�]�j h8��y���j��  Y�e� 3�@9����   ����E����} ��   �5 ��5<`�֋؉]Ѕ�th�5���֋��}ԉ]܉}؃��}�;�rK����9t�;�r>�7�֋���������5 ��֋��5����9]�u9E�t�]܉]ЉE؋��}ԋ]���E�a�}�as�E� ��t�ЃE����E�a�}�as�E�� ��t�ЃE����E������    �} u)���   j�  Y�u�����} tj��   Y�����Ë�U��j j�u������]�jj j ������Ë�U����3  �u�2  Yh�   ����̋�VW3�����<���u�����8h�  �0����`��tF��$|�3�@_^Ã$��� 3����S�,`V���W�>��t�~tW��W�`����& Y������|ܾ��_���t	�~uP�Ӄ�����|�^[Ë�U��E�4����4`]�jhX��>���3�G�}�3�9��u��2  j�+1  h�   �{���YY�u�4���9t���mj����Y��;�u�q����    3��Pj
�X   Y�]�9u+h�  W��`��uW菞��Y�<����    �]���>�W�t���Y�E������	   �E�������j
�)���YË�U��EV�4����> uP�#���Y��uj�A���Y�6�0`^]Ë�U���  ��  ���3ŉE��EV�uW3���4�����8�����0���9}u3��  ;�u�����8�����    �'�������  ������S�� �������L8$�����$�����?�����t��u'�M����u�@����  �%����    ������  �D8 tjj j V�  ��V蕑  Y����  ��D���  �����@l3�9H�� �����P��4����`3�;��`  ;�t8�?����P  ��`��4����� ���3���,���9E�#  ��@�����?������g  ���$���3���
��������ǃx8 t�P4�U�M��`8 j�E�P�K��P�ے  Y��t:��4���+�M3�@;���  j��D���SP�_�  �������  C��@����jS��D���P�;�  ������n  3�PPj�M�Qj��D���QP�� ���C��@����``�����=  j ��,���PV�E�P��$���� �4��`���
  ��@�����0������8���9�,�����  ����� ��   j ��,���Pj�E�P��$���� �E��4��`����  ��,�����  ��0�����8����   <t<u!�33Ƀ�
������@�����D��������<t<uR��D����̏  Yf;�D����I  ��8�������� t)jXP��D���蟏  Yf;�D����  ��8�����0����E9�@���������  ����8����T4��D8��  3ɋ�D8���  ��?��� ��D�����   ��4���9M��  ��3�+�4�����H���;Ms&�CA�� �����
u��0���� @F�@F���  rՋ���H���+�j ��(���PV��H���P��$���� �4��`���C  ��(����8���;��;  ��+�4���;E�l����%  ��?�����   ��4���9M�H  ��@��� ��+�4���j��H���^;MsC��Ή� �����
u�0���j[f��� �����@����@���f�Ɓ�@����  r�����H���+�j ��(���PV��H���P��$���� �4��`���i  ��(����8���;��a  ��+�4���;E�G����K  ��4�����,���9M�u  ��,�����@��� +�4���j��H���^;Ms;��,�����,���΃�
uj[f���@����@���f�Ɓ�@����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �``��;���   j ��(���P��+�P��5����P��$���� �4��`��t�(���;����@`��D���;�\��,���+�4�����8���;E�����?Q��(���Q�u��4����48��`��t��(�����D��� ��8�����@`��D�����8��� ul��D��� t-j^9�D���u�F���� 	   �N����0�?��D����R���Y�1��$���� �D@t��4����8u3��$�����    �����  ������8���+�0���[�M�_3�^�$�����jhx��L����]���u������  ����� 	   ����   ��x;�r�����  ����� 	   �3����ҋ����<� ��������D0��t�S苎  Y�e� ��D0t�u�uS�n������E���6���� 	   �>����  �M���E������   �E������Ë]S�ӎ  Y�jh���x����]���u������ 	   ����   ��x;�r������ 	   �o����ڋ����<� ��������D��t�S�Ǎ  Y�e� ��Dt1S�J�  YP��`��u�@`�E���e� �}� t�r����M��U���� 	   �M���E������   �E������Ë]S���  YË�U��V�u�F��t�t�v�\����f����3�Y��F�F^]�����w�����U��V������d����EtV����Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR����YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =RCC�t=MOC�t=csm�u*�������    �  �������    ~��������   3�]�jh�������}�]��   �s��s�u���������   �e� ;utb���~;w|��  �ƋO�4��u��E�   �|� t�sh  S�O�t��"  �e� ��u��+���YËe�e� �}�]�u��u���E������   ;ut�  �s�$���Ë]�u��(������    ~�������   Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�����3�A��  ���3��jh��m����M��t*�9csm�u"�A��t�@��t�e� P�q蕛���E������|����3�8E��Ëe��
  ̋�U��M�V�uƃy |�Q�I�42���^]Ë�U��3���;�u
�
  �A
  �E��E�9~OS�E�V�E�@�@��p� �M�q�P�GE�P�g�������u
K�������E��E�E�E�;|�^[�E���j��R�b�����������    t�
  �e� ��	  �M���	  �����Mj j ���   �D����j,hX��0����ً}�u�]�e� �G��E��v�E�P����YY�E��Z������   �E��L������   �E��>������   �3����M���   �e� 3�@�E�E��u�uS�uW�\������E�e� �o�E������Ëe��������   �u�}�~�   �O��O�^�e� �E�;Fsk��T;�~A;L;�F�L�QVj W�������e� �e� �u�E������E    �   �E��g�����E�맋}�u�E܉G��u��Z���Y�W����Mԉ��   �I����MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v�ܛ��Y��t�uV�*���YY�jh������3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w�O�  YY����   SV�>�  YY����   �G��M��QP�����YY���   �}�E�p�tH��  YY����   SV���  YY����   �w�E�pV谆�������   ���t|��W�9Wu8躉  YY��taSV證  YY��tT�w��W�E�p�d���YYPV�_������9肉  YY��t)SV�u�  YY��t�w�g�  Y��t�j X��@�E����  �E������E��3�@Ëe��  3��g����jh�������E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS������FP�w����YYP�vS������E�����������3�@Ëe���  ̋�U��} t�uSV�u�V������}  �uuV��u 蹖���7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP�C���]Ë�U���V�u�>  ���   W�X������    tG�J������   ����9t3�=MOC�t*=RCC�t#�u$�u �u�u�u�uV�Ԗ��������   �}� u�O  �u�E�P�E�PV�u W�����M���;M�sg���E�S�x�;7|G;p�B���H�Q��t�z u-�Y��@u%�u$�u�u j �u�u�u�u�����u�E����E��M����E�;M�r�[_^�Ë�U���4�MS�]�CVW�E� =�   �I��I�M����|;�|�  �u�csm�9>��  �~� ��)  �F;�t=!�t="��  �~ �  ��������    ��  ��������   �u��������   jV�E�v�  YY��u�  9>u&�~u �F;�t=!�t="�u�~ u��  �������    ��   �r������   �g����u3����   ����Y��u\3�9~�G�Lh���m~����uF��;7|��3  j�u�R���YY�EP�M��E���b���h���E�P�E̐�訋���u�csm�9>��  �~��  �F;�t=!�t="���  �}� ��   �E�P�E�P�u��u W�ٕ���M���;M���   �x�}�M��G��E�9��   ;O���   ��E�G��E��~r�F�@�X� �E��~#�v�P�u�E���������u�M��9E���M�E��}� ��.�u$�}��u �]��u��E��u�u�uV�u�����u�}���E��E����}�;E��P����}�} t
jV�����YY�}� ��   �%���=!���   �����   V�M���Y����   ���������������   �z����}$ �M���   Vu�u��u$�a����uj�V�u�u�]������v�g����]�{ v&�} ������u$�u �u�S�u�u�uV������ �������    t�T  _^[�Ë�U��V�u�����������^]� ��U��SVW�������   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������ 3�@_^[]�jh������������@x��t�e� ���3�@Ëe��E������λ������������@|��t������jh��J����5��<`��t�e� ���3�@Ëe��E������}����h�z�8`����������������U���SQ�E���E��EU�u�M�m��	�  VW��_^��]�MU���   u�   Q��  ]Y[�� ��U��   �em  ���3ŉE�SV�uWV�b�����3�Y������9F}�FjPPS��  ������������������|��s
������  ������ ���������� ��ÊH$����F  ������u�F�������+�ʋǋ��  ��V��+~���������[  �������  3�9P0�  �����9Vu�������������<  R�p,�p(�������+  ��������� ����;t(�3���;|,�)���j ������Qh   ������Q�4��`������j ��������������������  ����������������������������;��������������t7������K;�s+���u�J�;�s�H�9
u�������P��@��uЍ�����+�3����K  �@�t�V��:
u������B;�r������������u�������  ��x������    �%����F��   �V��u!�������   +N�@��<
��   jj j ��������  ��;�����u$;�����u�F�8��8
uG@;�r��F    �Yj �������������������  �����������������   ;�w�N��t
����   t�~������� �DtG������u��)����������� ������uѭ����������3������������M�_^3�[�6z����jh8��^���3�9E����u������    �p���������.�u虈��Y�e� �u�r���Y�E��U��E������   �E��U��M�����u�؈��YË�U��QQ�EV�u�E��EWV�E��${  ���Y;�u�R���� 	   �ǋ��J�u�M�Q�u�P��`�E�;�u�@`��t	P�D���Y�ϋ����� ������D0� ��E��U�_^��jhX��l�������]܉]��E���u������  ������ 	   �Ë��   ��x;�r������  ����� 	   �I����ы����<� ���������L1��t�P�z  Y�e� ��D0t�u�u�u�u��������E܉U���D���� 	   �L����  �]܉]��E������   �E܋U��������u��z  YË�U��V�uWV��y  Y���tP� ���u	���   u��u�@Dtj�y  j���y  YY;�tV�y  YP� `��u
�@`���3�V��x  ������ �����Y�D0 ��tW����Y����3�_^]�jhx�������]���u�l����  �Q���� 	   ����   ��x;�r�E����  �*���� 	   ������ҋ����<� ��������D0��t�S�%y  Y�e� ��D0tS�����Y�E�������� 	   �M���E������   �E�����Ë]S�}y  YË�U��9EuF�jP;Mu+�ݣ��YY���u3�]ËE�    �6�u�7�|�����Q�K�������tՉ�&3�@]Ë�U���EP�'������EYu��߃�]��Jx	�
�A�
�R����YË�U��S�U�������؃��t��P����Y��u��[]Ë�U���   ���3ŉE��M�EV�uW3��������|�����\�����P���ǅ$���^  ��0����������l���;�u�����    �;�������  ;�t��@@SurP�����Y������t���t�ȃ�������� �����A$u&���t���t�ȃ������ �����@$�t�����    ��������  �u������Ar���ƅ[��� ��t�����4�������  ����P趝��Y��t?��\�����t�����t�������Y���t��\���P�g���YYG�P�|���Y��u���  �<%�k  8G�X  3��������/�����T�����H�����d�����X�����Y�����c�����s�����Z�����k���ƅ{�����(���3�G���P�����Y��t��d�����H���k�
�DЉ�d�����   ��N��   ��   ��*tp��F��   ��It��Lut��{����   �O��6u�G�84u��(�������8�����<����m��3u�G�82u���\��dtW��itR��otM��xtH��Xu�A��c����9��ht(��lt��wt��s����"�G�8lt���{�����k������{�����k�����s��� �������c��� ��D���u������0�� �����������3���k��� ��@���ƅs��� u�<Stƅk����<Cuƅk������ ��L�����ntJ��ct��{t��\�����t�������Y���\�����t����W�����l�������  ��@�����D�����H�����t��d��� ��  ��o��  �_  ��c�  jdX;��K  ��  ��g~G��it!��n�{  ��c��� ��t�����
  ��
  ��L�����l�����-��  ƅY����  3ۃ�l���-u��P���� -C�	��l���+u��d�����\�����t����y�����l�����H��� u��d������l����k��d�����d�����tf��l�����P�����T������0���P��|���PCS��P�����$�������������
  ��\�����t����������l�����P�����Y��u���������   � � ��X���:�l�����   ��d�����d�������   ��\�����t���������P�����l�����X������0���P��|���PCS��P�����$�������������0
  ��l����k��d�����d�����tf��P�����l�����T������0���P��|���PCS��P�����$�������������	  ��\�����t����������l�����P�����Y��u���T��� �_  ��l���et��l���E�I  ��d�����d������5  ��P����e��0���P��|���PCS��P�����$������������D	  ��\�����t����_�����l�����-u,��P����-��0���P��|���PCS����������  �	��l���+u/��d�����d�����u!�d������\�����t����������l�����l����k��d�����d�����tf��P�����l�����T������0���P��|���PCS��P�����$����*��������j  ��\�����t���������l�����P茖��Y��u���t�����l����t��\�����l����K{��YY��T��� �  ��c��� �4  ��P�����4��������QP��@���� ��{���HP�5|��<`�Ѓ���  ��u��d���ǅH���   ��k��� ~ƅZ�����t�����l������t��\�����l����z��YY��H��� t��d�����d�������  ��\�����t���������l�������Q  ��ctL��su��	|	���9  �� u4��{�+  ��X���3ҋȃ�B������L�3ˋ�L������   ��c��� ��  ��Z��� ��  �� �����P��m  Y��t��\�����t����������!��������P�����ǅ���?   ���   �� ���P�����P�'l  f�������f����e  �Ã�p��  �������HH��  ���������t3�;�l�����  ��[�����c��� �K  �� ���������:  ��k��� ~ƅZ����^�wu
�wƅX����j �E�j P�l�����>]u�]F�E� �   ��/����   F<-uq��tm���]tfF:�s��{������{�����:�{���s,��{���*����Ћσ��ǳ�����D�GJu苝L�����{�������������D�2���ȊЋ���������D���L����<]�c������  ��D�����@����b�����+u.��d���u��t	ƅs������\�����t��������؉�l�����0��  ��\�����t���������؉�l�����xt_��XtZ��L���xǅT���   t&��H��� t��d���u��s���ǅL���o   �.  ��t������t��\���S�w��YYj0[�  ��\�����t����l�����H��� �؉�l���t��d�����d���}��s���ǅL���x   ��   �F��@����x���G�r�����t������t��\���P�w��YY;���  ��c��� ��  ��4�����c��  ��Z��� t��@���3�f���  ��@����  �  ƅ{�����l�����-u	ƅY������+u.��d���u��t	ƅs������\�����t����x����؉�l�����(��� �<  ��s��� ��   ��L���xt]��L���ptT��P�Q���Y����   ��L���ou��8��   ��8�����<��������Kj j
��<�����8����o  �����0��P聑��Y��tk��8�����<�����S��������Y��l�����T����CЙ����H��� ��8�����<���t��d���t7��\�����t��������؉�l����!�����t������t��\���S�Zu��YY��Y��� �������   ��8�����<����؃� �ى�8�����<�����   ��s��� �������   ��L���xt/��L���pt&��P����Y��tq��L���ou
��8}c���%k�
� ��P�m���Y��tKS��������Y��l�����T�����H��� �|�t��d���t7��\�����t��������؉�l����o�����t������t��\���S�ft��YY��Y��� t�߃�L���Fu��T��� ��T��� �  ��c��� u8��4�����@�����(��� t��8������<����F���{��� t�>�f�>��D�����[���G��D����d<%u8GuG��\�����t�����������G��l�����D���;�uw��P�g  Y��t%��\�����t��������G��D���;�u7��t�����l����u�?%uN��D����xnuB�����������4��l��������t��\���P�@s��YY���t��\�����l����(s��YY��0���u��P����p��Y��l����u*��4�����u8�[���u�������� t%������ap������� t
������`p���4���[�M�_3�^�?f���Ë�U���V�u�M��&c���E�u��t�0��u$�ʶ���    �m����}� t�E�`p�3���  �} t�}|Ѓ}$ʃe� �M�S�W�~���   ~�E�P��jP��  �M������   ���B����t�G�ǀ�-u�M���+u�G�E���O  ���F  ��$�=  ��u*��0t	�E
   �6�<xt<Xt	�E   �#�E   �
��u��0u�<xt<Xu�_�����3��u���   �U����N�у�t�˃�0���  t0�K�����w�� ���;Ms�M9E�r(u;M�v!�M�} u#�EO�u �} t�}�e� �[�U��UщU��G늾����u�u=��t	�}�   �w	��u+9u�v&�*����E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�_[^�Ë�U��3�P�u�u�u9,�uh���P������]Ë�U��3��M;�(�t
@��r�3�]Ë�,�]Ë�U����  ���3ŉE�SV�uWV������3�Y�����;��l  j�m  Y���  j�m  Y��u�=$���   ���   �6  hd�h  � �W�vl  ������   h  �R�VSf�Z���`��  ��uh4�SV�>l  ����t3�PPPPP�	���V�
l  @Y��<v*V��k  �E����+�j��h,�+�SP�k  ����u�h$��  VW�j  ����u������VW�rj  ����u�h  h؋W��h  ���^SSSSS�y���j���`��;�tF���tA3��G�����f9Gt@=�  r�S�����P�����P�]�����YP�����PV��`�M�_^3�[�b����j�k  Y��tj�k  Y��u�=$�uh�   �%���h�   ����YYË�U���   ���3ŉE��}�ESVW�}��x�����   ��t��� h�   ��|�����Q�u�uP�:l  ������ub�@`��zuxVV�u�u��x����l  ����p�����tXFVP�N�����YY��tH��p�����t���S�u�u��x�����k  ������tjV�����3�YY;�u!9�t���tS�k��Y����M�_^3�[��`���ÍN�QSVP��(  ����u9�t���tS��j��Y3���WWWWW�ΰ���}uH�5�`3�PP�u��u�֋؅�tjS蔍��YY���tSP�u�u�օ�u��7�zj���' Y�p����} �f�����x��� j��x���P�E    P�u��`���<�����x�����c�����U��E�H�]Ã=� u蔦��V�5�W3���u����   <=tGV襚��Y�t���u�jGW�ی����YY�=����tˋ5�S�3V�t����>=Y�Xt"jS譌��YY���t?VSP�>_������uG���> u��5��i���%� �' ���   3�Y[_^��5���^i���%�� �����3�PPPPP�U���̋�U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�%j  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�@i  Y��t��M�E�F��M��E���i  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9�u����h  �P�VS�T���`�$��5��;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�������Y;�t)�U��E�P�WV�}�������E���H����5��3�����_^[�Ë�U���SV��`��3�;�u3��wf93t��f90u���f90u�W�=``VVV+�V��@PSVV�E��׉E�;�t8P�Q���Y�E�;�t*VV�u�P�u�SVV�ׅ�u�u��wf��Y�u�S��`�E��	S��`3�_^[�Ë�V�t��t�W��;�s���t�Ѓ�;�r�_^Ë�V�|��|�W��;�s���t�Ѓ�;�r�_^Ë�U��V���������2  �N\�U��W9t�����   ;�r���   ;�s9t3���t�P��u3���   ��u�` 3�@��   ����   �MS�^`�N`�H����   j$Y�~\�d9 �����   |� �~d=�  �u	�Fd�   �~=�  �u	�Fd�   �n=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=� �u	�Fd�   �=� �u�Fd�   �vdj��Y�~d��` Q��Y�^`[���_^]Ë�U��csm�9Eu�uP����YY]�3�]Ë�U�������e� �e� SW�N�@��  ��;�t��t	�У���eV�E�P�a�u�3u��a3��T`3�� a3��E�P��`�E�3E�3�;�u�O�@����u��G  ����5���։5��^_[�Ë�U��E�X�]Ë�U���5X��<`��t�u��Y��t3�@]�3�]Ë�U���(3��E��E�9`�t�5���<`�����M��   V;���  ��  ���  �  jZ+���   I��   ����   I��   ����   ItN��	�  �E�   �E���M��M�u�]���M��]�Q��]���Y����  �©��� "   ��  �E����M��M�u�]���M��]�Q��E�   �]���Y�  �E�   �E�����E���M�u��M�]���]���?  �U��E���W����E���ΉU��E���?����E���q�����tWItHIt9It ��t���  �E�܍��E�ԍ��E���M��u��u����E���c����E�   �������E���   �E�   �E�̍�������������   �$���E����E����E�����E�č��Eܼ��t����Eܴ��h����Eܬ��\����Eܨ���Eܤ���Eܠ��M��u�M����M�]���]�M��]�Q�E�   ��Y��u������ !   �E��^�Ðp�y���������#����������ʡj
��`���3�Ë�U��QQSV���  V�5��j  �EYY�M�ظ�  #�QQ�$f;�uU�Pi  YY��~-��~��u#�ESQQ�$j��g  ���tVS�nj  �EYY�f�ES��d���\$�E�$jj�A�h  �]��E�Y�EY������DzVS�*j  �E�YY�"�� u��E�S���\$�E�$jj�g  ��^[�Ë�U��� �e� Wj3�Y�}��9Eu详���    �R�������x�MV�u��t��u苦���    �.�������S�����E�;�w�M��u�E��u�E�B   �u�u�P�u��k  ������t�M�x�E��  ��E�Pj 蛺��YY��^_�Ë�U���uj �u�u�u�<�����]Ë�U��} u������    蚥�����]��uj �5���a]�����U���0���S�ٽ\�����=`� t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=`� t�#  ��8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8����3  �   [�À�8�����=� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   ������������������s4�(��,ǅr���   ������������� �����v� �VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�t  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����K   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[��������̀zuf��\���������?�f�?f��^���٭^����L��剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����L��剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����D����۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-0���p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR��q  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��`��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z���������������|������   s�������������������t������   v����떋�U���S�u�M���K���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�N  YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�  �� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U��QQ���3ŉE�S3�VW�]�9]u�E� �@�E�5h`3�9] SS�u���u��   P�u�֋�;�u3��~<�����w4�D?=   w輞����;�t� ��  �P��l��Y;�t	� ��  ���؅�t��?Pj S�M����WS�u�uj�u�օ�t�uPS�u�a�E�S�2J���E�Y�e�_^[�M�3��AM���Ë�U����u�M��)J���u$�E��u�u�u�u�uP��������}� t�M��ap��Ë�U��M��tj�3�X��;Es蘝���    3�]��MV���uF3����wVj�5���\`��u2�=\� tV����Y��uҋE��t�    3���M��t�   ^]Ë�U��} u�u�k��Y]�V�u��u�u�ZV��Y3��MW�0��uFV�uj �5���a����u^9\�t@V�.���Y��t���v�V����Y�Ĝ���    3�_^]�賜�����@`P�c���Y���蛜�����@`P�K���Y����ʋ�U��MS3�;�vj�3�X��;Es�f����    3��A�MVW��9]t�u�@���Y��V�u������YY��t;�s+�Vj �S�K������_^[]Ë�U���S�XBV���HD�M���u�����  �e� W�E�FPj1S�E�jP�L������FPj2S�E�jP�8�����FPj3S�E�jP�$�����FPj4S�E�jP������P��FPj5S�E�jP�������FPj6S�E�jP�����Vj7S��E�jP�������F Pj*S�E�jP�������P��F$Pj+Sj�E�P������F(Pj,S�E�jP������F,Pj-S�E�jP������F0Pj.S�E�jP�m�����P��F4Pj/S�E�jP�V�����FPj0S�E�jP�B�����F8PjDS�E�jP�.�����F<PjES�E�jP������P��F@PjFS�E�jP������FDPjGS�E�jP�������FHPjHS�E�jP�������FLPjIS�E�jP�������P��FPPjJS�E�jP������FTPjKS�E�jP������FXPjLS�E�jP������F\PjMS�E�jP�t�����P��F`PjNS�E�jP�]�����FdPjOS�E�jP�I�����FhPj8S�E�jP�5�����FlPj9S�E�jP�!�����P��FpPj:S�E�jP�
�����FtPj;S�E�jP�������FxPj<S�E�jP�������F|Pj=S�E�jP�������P����   Pj>S�E�jP��������   Pj?S�E�jP��������   Pj@S�E�jP��������   PjAS�E�jP�o�����P����   PjBS�E�jP�U�������   PjCS�E�jP�>�������   Pj(S�E�jP�'�������   Pj)S�E�jP������P����   Pj�u��E�jP���������   Pj �u��E�jP���������   Ph  �u��E�jP��������   Ph	  �u��E�j P������E���P���   ���   Pj1S�E�jP��������   Pj2S�E�jP�i�������   Pj3S�E�jP�R�������   Pj4S�E�jP�;�����P����   Pj5S�E�jP�!�������   Pj6S�E�jP�
�������   Pj7S�E�jP���������   Pj*S�E�jP�������P����   Pj+S�E�jP���������   Pj,S�E�jP��������   Pj-S�E�jP��������   Pj.S�E�jP�}�����P����   Pj/S�E�jP�c�������   Pj0S�E�jP�L�������   PjDS�E�jP�5�������   PjES�E�jP������P����   PjFS�E�jP��������   PjGS�E�jP��������   PjHS�E�jP��������  PjIS�E�jP������P���  PjJS�E�jP�������  PjKS�E�jP�������  PjLS�E�jP�w������  PjMS�E�jP�`�����P���  PjNS�E�jP�F������  PjOSj�E�P�/������   Pj8S�E�jP�������$  Pj9S�E�jP������P���(  Pj:S�E�jP��������,  Pj;S�E�jP��������0  Pj<S�E�jP�������4  Pj=S�E�jP������P���8  Pj>S�E�jP�������<  Pj?S�E�jP�q������@  Pj@S�E�jP�Z������D  PjAS�E�jP�C�����P���H  PjBS�E�jP�)������L  PjCS�E�jP�������P  Pj(S�E�jP��������T  Pj)Sj[�E�SP�������P���X  Pj�u��E�SP��������\  Pj �u��E�SP������`  Vh  �u���E�SP������<�_^[�Ë�U��V�u���c  �v�MM���v�EM���v�=M���v�5M���v�-M���v�%M���6�M���v �M���v$�M���v(�M���v,��L���v0��L���v4��L���v��L���v8��L���v<��L����@�v@��L���vD��L���vH�L���vL�L���vP�L���vT�L���vX�L���v\�L���v`�L���vd�L���vh�{L���vl�sL���vp�kL���vt�cL���vx�[L���v|�SL����@���   �EL�����   �:L�����   �/L�����   �$L�����   �L�����   �L�����   �L�����   ��K�����   ��K�����   ��K�����   ��K�����   ��K�����   ��K�����   �K�����   �K�����   �K����@���   �K�����   �K�����   �|K�����   �qK�����   �fK�����   �[K�����   �PK�����   �EK�����   �:K�����   �/K�����   �$K�����   �K�����   �K����   �K����  ��J����  ��J����@��  ��J����  ��J����  ��J����  �J����  �J����   �J����$  �J����(  �J����,  �J����0  �|J����4  �qJ����8  �fJ����<  �[J����@  �PJ����D  �EJ����H  �:J����@��L  �,J����P  �!J����T  �J����X  �J����\  � J����`  ��I����^]Ë�U��SV�u�~  W���tBhd  j��l����YY��u3�@�I�Ƌ��R�����tW�G���W�I��YY��Ǉ�      ������   ;�t�   P� `���   3�_^[]Ë�U��V�u��tY�;8�tP�UI��Y�F;<�tP�CI��Y�F;@�tP�1I��Y�F0;h�tP�I��Y�v4;5l�tV�I��Y^]Ë�U���SV�uW3��u��}�9~u9~u�}��}��8��e  jPj��k����YY;�u3�@�  ���   jY��j��dk��3�Y�E�;�u	S�H��Y�ыu�89~��   j�<k��Y�E�;�u3�FS�sH���u��kH��YY���D  �8�v>SjV�E�jP�q������CPjV�E�jP�]�����CPjV�E�jP�I�����C0PjV�E�jP�5�����P��C4PjV�E�jP�������tS�{���Y����k����C����0|��9��0�@�8 u��>��;u���N�F�> u���8���<��C�@��C�h��C0�l��}��C4�M��u3�@��M���t����   �= `��tP�׋��   ��tP�ׅ�u���   �EG�����   �:G��YY�E����   �E����   ���   3�_^[�Ë�U��V�u����   �F;D�tP��F��Y�F;H�tP��F��Y�F;L�tP��F��Y�F;P�tP��F��Y�F;T�tP�F��Y�F ;X�tP�F��Y�F$;\�tP�F��Y�F8;p�tP�yF��Y�F<;t�tP�gF��Y�F@;x�tP�UF��Y�FD;|�tP�CF��Y�FH;��tP�1F��Y�vL;5��tV�F��Y^]Ë�U���SV�uW3��}��u��}�9~u9~u�}��}��8���  jPj��h����YY;�u3�@�  j�h��Y�E�;�u	S�E��Y���89~�4  j�]h��Y�E�;�uS�E���u��E��Y�҉8�v8�CPjV�E�jP�������CPjV�E�jP������CPjV�E�jP�p�����CPjV�E�jP�\�����P��CPjV�E�jP�E�����C PjPV�E�jP�1�����C$PjQV�E�jP������C(PjV�E�j P�	�����P��C)PjVj �E�P�������C*PjTV�E�j P�������C+PjUV�E�j P�������C,PjVV�E�j P������P��C-PjWV�E�j P������C.PjRV�E�j P������C/PjSV�E�j P�w�����C8PjV�E�jP�c�����P��C<PjV�E�jP�L�����C@PjV�E�jP�8�����CDPjV�E�jP�$�����CHPjPV�E�jP������P��CLPjQV�E�jP��������t$S����S��C���u��C���u��C����������C����0|��9��0�@�8 u�� ��;u���N�F�> u���jY�8����E���   �	����   �I�u�K���   �I�K���   �I0�K0���   �@4�M��C43�@3��9}�t�M�����   ;�tP� `���   ;�t#P� `��u���   ��B�����   ��B��YY�E����   �E����   ���   3�_^[��3�Ë�U��MVW��t�}��u�Q���j^�0��������A�U��u� ���> tFOu���t�+��B��tOu��u� ����j"Y����3�_^]���������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^�Ë�U��ES3�VW9]u;�u9]u3�_^[]�;�t�};�w�x���j^�0��������9]u��ҋU;�u��ك}���u��+�
�B:�t"Ou����+���A:�tOt�Mu�9]u�;�u��}�u�MjP�\�X�x���������j"Y���낋�U��3�S3�@9]|FVW��t>�EÙ+��E���<��7�E�0�Z  YY��u
�M���9�yN�u��^;]~�_^3Ʌ���[��]Ë�U��Q��tP�> tKh��V��u��YY��t:h��V��u��YY��uj�E�Ph   �w��`��t)�E���V�S��Y�E���j�E�Ph  �w��`��u3��Ã}� u��p`�Ë�U��3�f�Mf;�p�t����r�3�@]�3�]Ë�V3�� �A�B<w����
�A�<w�������t�Њ
��uڋ�^�3��
B��A|��Z~��a��w@��Ë�U���|���3ŉE�VW�}�W����׋�������jx�E�P���   ���%���  PW�a��u	!��   @�A�E�P���   �0Y  YY��uW����Y��t���   ���   ���   ���   ���Ѓ��M�_3�^�E5���� ��U��QV��j�E�P��%�  h      P��`��u3��);u�t!�} t�E�0W�������V���o��Y;�_t�3�@^�Ë�U���|���3ŉE�SVW�}�T����׍��   �����a��jx�E�P�F���%���  PW�Ӆ�u�f 3�@�c  �E�P�v�*X  YY����   jx�E�P�F���%���  PW�Ӆ�t��E�P�6��W  YY��u�N  �~�R�FuO�F��t,P�E�P�6��X  ����u�6�N�~�n��Y;Fu!�~��V��uW����Y��t	���V�~�N�   #�;���   jx�E�P�F���%���  PW�Ӆ������E�P�6�OW  Y3�Y��u0�N   �F9^t
   �F�H9^t<�6�+n��Y;Fu/Vj�9^u49^t/�E�P�6�W  YY��uVS������YY��t�N   9^u�~�F���Ѓ��M�_^3�[�3���� ��U���|���3ŉE�VW�}�~���׍��   ������jx�E�P�F���%���  PW�a��u!F@�\�E�P�6�cV  YY��u
9Fu1Vj��~ u0�~ t*�E�P�6�<V  YY��uVP���?���YY��t
�N�~�~�F���Ѓ��M�_3�^�Y2���� �6�m���v�����@�F��l��������f @�~ YY�FtjX������jhd��F� a�F�   t�   t�u�f ��6�l�������@Y�FtjX�������jh5��F� a�Fu�f Ë�U��SVW�0}�����   �E��u�O  ��   ���@�_�t�8 tSjh���/�������g ��t[�8 tV���t�8 t	�����������S���� ��   Wj@h�����������tf���t�; t	�������R�������I���t0�; t+S�k������Y�j@hb��G� a�Gu�g ��G  �a�G�G� ��   �u�ƃ����#���������u����   ����  ��   ����  ��   ��P�x`����   j�w�$a����   �E��tf�Of�f�Of�Hf�p�]��th�5a�  f9u h��j@S�/������t3�PPPPP����j@Sh  �w�օ�t,j@�C@Ph  �w�օ�tj
j��S�u�U  ��3�@�3�_^[]Ë�U��VW�}�ǃ� ��  H��  H�l  H�!  H��  �M�ESj Z�2  �0;1tt�0�+�t3ۅ��Ít����+  �p�Y+�t3ۅ��Ít����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít��3�����  �p;qtv�p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít����e  �p�Y+�t3ۅ��Ít��3����B  �p;qtv�p�Y+�t3ۅ��Ít����  �p	�Y	+�t3ۅ��Ít�����  �p
�Y
+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít��3�����  �p;qtv�p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít����t  �p�Y+�t3ۅ��Ít����U  �p�Y+�t3ۅ��Ít��3����2  �p;qtv�Y�p+�t3ۅ��Ít����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít��3�����  �p;qtv�p�Y+�t3ۅ��Ít�����  �p�Y+�t3ۅ��Ít����d  �p�Y+�t3ۅ��Ít����E  �p�Y+�t3ۅ��Ít��3����"  �p;qtv�p�Y+�t3ۅ��Ít�����   �p�Y+�t3ۅ��Ít�����   �p�Y+�t3ۅ��Ít�����   �p�Y+�t3ۅ��Ít��3�����   �p;qtj�p�Y+�t3ۅ��Ít���uw�p�Y+�t3ۅ��Ít���u\�p�Y+�t3ۅ��Ít���uA�p�Y+�t3ۅ��Ít��3���u"��+�;�������σ���  �$�]����  �P�;Q�ti���Q�+�t3҅��t���u��p��Q�+�t3҅��t���u��p��Q�+�t3҅��t���u��p��Q�+�t3҅��t��3���u��P�;Q�tu���Q�+�t3҅��t����\����p��Q�+�t3҅��t����=����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����t����P�;Q�tu���Q�+�t3҅��t����N����p��Q�+�t3҅��t����/����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����e����P�;Q�tu���Q�+�t3҅��t����?����p��Q�+�t3҅��t���� ����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tm���Q�+�t3҅��T���u6�p��Q�+�t3҅��T���u�p��Q�+�t3҅��T���t����@��I�+�t3Ʌ����D	��3���u3�[�  �P�;Q�tu���Q�+�t3҅��t����5����p��Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t����p����p��Q�+�t3҅��t��3����M����P�;Q�tu���Q�+�t3҅��t����'����p��Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t����b����p��Q�+�t3҅��t��3����?����P�;Q�tu���Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t���������p��Q�+�t3҅��t����r����p��Q�+�t3҅��t����S����p��Q�+�t3҅��t��3����0����P�;Q�tu���Q�+�t3҅��t����
����p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������I��@�+��8���3Ʌ����D	��(����P�;Q�tu���Q�+�t3҅��t����c����p��Q�+�t3҅��t����D����p��Q�+�t3҅��t����%����p��Q�+�t3҅��t��3��������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����{����P�;Q�tu���Q�+�t3҅��t����U����p��Q�+�t3҅��t����6����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����m����P�;Q�tu���Q�+�t3҅��t����G����p��Q�+�t3҅��t����(����p��Q�+�t3҅��t����	����p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t���������Q��p�+�t3҅��t���������Q��p�+�t3҅��t���������Q��p�+�t3҅��t��3����^����P�;Q�tu���Q�+�t3҅��t����8����p��Q�+�t3҅��t��������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3��������f�P�f;Q��f����Q��p�+�����3҅��T�����  ������P�;Q�tv�Q��p�+�t3҅��t����z����p��Q�+�t3҅��t����[����p��Q�+�t3҅��t����<����p��Q�+�t3҅��t��3��������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t����l����p��Q�+�t3҅��t����M����p��Q�+�t3҅��t����.����p��Q�+�t3҅��t��3��������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3���������P�;Q�tv�Q��p�+�t3҅��t����]����p��Q�+�t3҅��t����>����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������P�;Q�tu���Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t���������p��Q�+�t3҅��t��3����u����P�;Q�tu���Q�+�t3҅��t����O����p��Q�+�t3҅��t����0����p��Q�+�t3҅��t��������p��Q�+�t3҅��t��3���������p��Q�+�����3҅��T����������c����M�u��+�t3҅��D�����   �A�V+�t3҅��D�����   �A�V+�t3҅��D�����   �A�N+���   3Ʌ����D	��   �M�u��+�t3҅��D���ud�A�V+�t3҅��D���uI�A�N뤋M�u��+�t3҅��D���u �A�N�x����E�M� �	�g���3�_^]Ë���n�@�)�9���������_�1��*���������Q�#�����������C���������v����U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�ø@�ø��Ë�U������S3�V�u�E��]�]��]��F�> t��<at,<rt"<wt�j���    �<j��3��F  �  ��M��	�	  �M�3�AF�W����  �y� @  ���  ����S��   t�� ��   ��tRHtC��t-��
t!����  9E���   �E�   ����   ��   ��@��   ��@�   �E�   �   ����   �E���������ǉE��   �}� ut�E�   �� �n��TtZ��tEHt0��t���  �� �  uE��G�}� u;�e������E�   �1�}� u%	U��E�   ��� �  u�� �  ��   ��t3���F���������}� ��   �F�> t�jVhؙ��I  ����u~���F�> t��>=unF�> t�jhܙV�dH  ����u����   �?jh�V�EH  ����u����   � jh�V�&H  ����u����   �F�> t��> t�h���    �4h���h�  �u�ES�uP�E  ����t3��"���E�M��H3ɉH��H�H�M�H_^[��jh���z��3�3��}�j����Y�]�3��u�;5@
��   �(���9t[� �@��uH� �  uA�F���w�FP����Y����   �(��4�V��%��YY�(����@�tPV�H&��YYF둋��}��cj8�C��Y�(���;�tNh�  �(����� P��`���(�u�4�� ��Y�(�������� P�0`�(��<��}�_;�t�g �  �_�_��_�O��E������   ����y��Ë}�j�+���Y�����������SVW�T$�D$�L$URPQQh��d�5    ���3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�B  �   �C�T  �d�    ��_^[ËL$�A   �   t3�D$�H3����U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�  3�3�3�3�3���U��SVWj Rh6�Q�l  _^[]�U�l$RQ�t$������]� ��U��V�uV�d  Y���u�e��� 	   ����MW�uj �uP��`�����u�@`�3���tP�e��Y���������� ������D0� ���_^]�jh���w���]���u�3e���  �e��� 	   ����   ��x;�r�e���  ��d��� 	   �d���ҋ����<� ��������D0��t�S��  Y�e� ��D0t�u�uS��������E���d��� 	   �d���  �M���E������   �E��6w��Ë]S�4  YË�U���SW�}3�;�u�Md���    ��c������e  VW�v����Y�u�9_}�_jSV��������E�;���   �W��  u+G�%  ��O��+ى]���t<������ ������D2�t��;�s���:
uCB;�r��]�}� u����   ��x��c���    �   �G��   �W��u!U��   �]��u�+�������� ��E����D0�tyjj �u�������;E�u �G�M��	�8
u�E@;�r��G    �@j �u��u����������y����8�   9Ew�O��t��   t�G�E��D0t�E�E)E��E�E�^_[�Ë�U��E�l��p��t��x�]Ë�U��E�4�V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5t��<`�j hؾ��t��3��}�}؋]��Kt��jY+�t"+�t+�tY+�uC�\�����}؅�u����T  �l��l��U�w\���]���Y�p��Q�Ã�t2��t!Ht��a���    �a��빾t��t���p��p��
�x��x��E�   P�<`�E�3��}���   9E�uj��z��9E�tP�|��Y3��E���t
��t��u�O`�MԉG`��u>�Od�M��Gd�   ��u,�(��M܋,�(�9M�}�M�k��W\�D�E����PZ����E������   ��u�wdS�U�Y��]�}؃}� tj �{��Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3��s��Ã%�� �����Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �������U��W�}3�������ك��E���8t3�����_�Ë�U���SV�u�M�����]�   ;�sT�M胹�   ~�E�PjS�����M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�<  YY��t�Ej�E��]��E� Y��_��� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�4����$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=,� u�E�H���w�� ]�j �u�����YY]Ë�U���(���3ŉE�SV�uW�u�}�M��C���E�P3�SSSSW�E�P�E�P�yJ  �E�E�VP��?  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�����Ë�U���(���3ŉE�SV�uW�u�}�M��
���E�P3�SSSSW�E�P�E�P��I  �E�E�VP�sD  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[����Ë�U��MS�YV�u3�;�u�]��j^�0�[]�����   9Ev�U�;�~��@9Ew�]��j"Y�����W�~�0�ǅ�~���t��C�j0Y�@J���M�  ��x�;5|�� 0H�89t�� �>1u�A�W�2G��@PWV�����3�_^[]Ë�U��Q�M�AS����% �  V��  #�W�E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��B��<  �U����������U��E����������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0���3ŉE��ES�]V�E�W�EP�E�P�"���YY�E�Pj j���uЋ���f��N  �u܉C�E��E��C�E�P�uV��
����$��u�M�_�s^��3�[�7����3�PPPPP�;[�����������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�*t��YË�U��E�M%����#�V�u������t$��tj j �4W  YY��Z��j^�0�8Z�����P�u��t	�W  ���W  YY3�^]Ë�U����UV�uj�X�E�U�;�u�[Z���  �@Z��� 	   ����}  S3�;�|;5�r�1Z����Z��� 	   �Y������N  ����W���<� �����L0��u��Y�����Y��� 	   �h�����wN�]�;��  ����  9]t5�D0$����E���HjYtHu���Шt����U�]�]��z���Шu�Y����pY���    �Y���6����M;�r�E�u�R5����Y�]���u�>Y���    �FY���    ����n  jj j �u蚎����D(���T,���AH��tz�I��
tr�} tl�M�}� ���C�E�   �D
tP��L%��
tE�} t?��@�M�}��E�   �D%
u%��L&��
t�} t��@�M�E�   �D&
j �M�Q�uP��4��`���x  �M���m  ;M�d  �M�D� ���  �}��  ��t
�;
u��� ��]��E�É]�E�;���   �M�<��   <t�CA�M�   �E�H;�s�A�8
u���M�
�u�E�m�Ej �E�Pj�E�P��4��`��u
�@`��uE�}� t?��DHt�}�
t����M��L�%;]�u�}�
t�jj�j��u�������}�
t�C�E�9E�F������D� @u����C��+E��}��E���   ����   K���xC�   3�@�����;]�rK�@��P� t�����P���u��V��� *   �zA;�u��@��D1Ht%C�T1��|	���T%C��u	���T&C+���ؙjRP�u�������E�+]���P�uS�u�j h��  �h`�E��u4�@`P�V��Y�M���E�;EtP���Y�E�����  �E��  �E�3�;�����E�L0�ƅ�tf�;
u��� ��]��E�É]�E�;��  �E�����   ��tf������E�   �M���;�s�Hf�9
u���Ej
�   �M�   �Ej �E�Pj�E�P��4��`��u
�@`��u[�}� tU��DHt(f�}�
t�jXf���M��L��M��L%��D&
�*;]�uf�}�
t�jj�j��u跊����f�}�
t	jXf����E�9E�������t�@u��	f� f���+]��]������@`j^;�u��T��� 	   ��T���0�j�����m�Z����e� �\���3�_[^��jh���&g���]���u�T���  �T��� 	   ����   ��x;�r�T���  �jT��� 	   �T���ҋ����<� ��������D0��tƸ���;E�@u�>T���  �#T���    �S�C  Y�e� ��D0t�u�uS�������E����S��� 	   ��S���  �M���E������   �E��f��Ë]S�  Y������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��t�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h�h�\d�    P��SVW���1E�3�P�E�d�    �e��E�    h   �*�������tT�E-   Ph   �P�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE�3ҁ9  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U��E���u�RR��� 	   3�]Å�x;�r�7R��� 	   ��Q���ދȃ����� ����D��@]Ë�U��E���]Ë�U��Q�=���u�Q  ������u���  ��j �M�Qj�MQP�,a��t�f�E�Ë�U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M�������E�9Xu�E;�t�f�8]�t�E��`p�3�@�ˍE�P�P��   YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�h`���E�u�M;��   r 8^t���   8]��f����M��ap��Z�����P��� *   8]�t�E��`p�����;���3�9]��P�u�E�jVj	�p�h`���:���뺋�U��j �u�u�u�������]Ë�U����u�M�������E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U��EVW��xY;�sQ���������<� �����<�u5�=$�S�]u�� tHtHuSj��Sj��Sj��0a��3�[���O��� 	   ��O���  ���_^]Ë�U��MS3�VW;�|[;�sS��������<� �����D0t6�<0�t0�=$�u+�tItIuSj��Sj��Sj��0a���3���PO��� 	   �XO������_^[]Ë�U��E���u�<O���  �!O��� 	   ���]Å�x;�r�O���  ��N��� 	   �N���Ջ����� ������Dt͋]�jh8��Fa���}����������4� ��E�   3�9^u5j
�i��Y�]�9^uh�  �FP��`��u�]��F�E������0   9]�t���������� ��D8P�0`�E��a���3ۋ}j
�Th��YË�U��E�ȃ����� ����DP�4`]�jhX��`���M��3��}�j�&h��Y��u����a  j��h��Y�}��}؃�@�;  �4� �����   �u��� �   ;���   �Fu[�~ u8j
�h��Y3�C�]��~ uh�  �FP��`��u�]���F�e� �(   �}� u�^S�0`�FtS�4`��@냋}؋u�j
�Rg��YÃ}� u��F��+4� ���������u�}��uyG�,���j@j �E)��YY�E���ta�� ���� ���   ;�s�@ ���@
�` ��@�E������}�����σ����� ��DW�����Y��u�M���E������	   �E��B_���j�f��YË�U��3�@�} u3�]��U��SVWUj j h���u�R  ]_^[��]ËL$�A   �   t2�D$�H�3��j���U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��d�5    ���3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ�P��SQ�P��L$�K�C�kUQPXY]Y[� �����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U���$���3ŉE��ES�E��EVW�E��JC���e� �=�� �E�u}h���(a�؅��  �=�`h��S�ׅ���   �58`P��h��S�����P��hx�S�����P��h\�S�����P�֣����thD�S��P�֣������M�5<`;�tG9��t?P���5�����֋؅�t,��t(�ׅ�t�M�Qj�M�QjP�Ӆ�t�E�u	�M    �3���;E�t)P�օ�t"�ЉE��t���;E�tP�օ�t�u��ЉE��5���օ�t�u�u��u��u����3��M�_^3�[�+����Ë�U��V�uW��t�}��u��H��j^�0�iH����_^]ËM��u3�f��݋�f�: t��Ou��t�+��f�
��f��tOu�3���u�f��sH��j"Y���몋�U��US�]VW��u��u9Uu3�_^[]Å�t�}��u�8H��j^�0��G�����݅�u3�f��ЋM��u3�f��ԋ��u��+��f���f��t'Ou��"��+��f���f��tOtKu��u3�f����y���3����u�MjPf�DJ�X�d���f��G��j"Y����j�����U��Ef���f��u�+E��H]Ë�U��V�uW��t�}��u�hG��j^�0�G����_^]ËE��uf��ߋ�+��f���f��tOu�3���u�f��(G��j"Y���뼋�U��M��x��~��u� �]á �� �]���F���    �F�����]Ë�U������3ŉE��E� �@SVW�=�`3�VV�u�E��u�׋ȉM�;�u3��   ~Ej�3�X���r9�D	=   w��F����;�t����  ���P���Y;�t	� ��  �����3�;�t��u�S�u�u�ׅ�t VV9uuVV��u�uj�SV�u��``��S�B���Y�ƍe�_^[�M�3��R����Ë�U����u�M��:����u�E��u�u�uP��������}� t�M��ap��Ë�U����u�M�� ����E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�c  �EPSj �u�H`�M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�  Y����  �t�Etj�y  Y����x  ����   �E��   j�W  �EY�   #�tT=   t7=   t;�ub��M����`���{L�H��M�����{,�`��2��M�����z�`����M�����z�P���P���������   ���   �E��   3��t��W�}���������D��   ��E�PQQ�$�  �M��]�� �����������}�E����c�S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj�   Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}�f@��� "   ]��Y@��� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���h�;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�I�������uV�,���Y�E�^�Ë�l��h��  �u(�  �u�����E ���Ë�U��=`� u(�u�E���\$���\$�E�$�uj�/�����$]��B?��h��  �u� !   �\  �EYY]Ë�S��QQ�����U�k�l$���   ���3ŉE��s �CP�s��������u#�e��P�CP�CP�s�C �sP�E�P�j������s�o������=`� u+��t'�s �C���\$���\$�C�$�sP�q�����$�P�����$��  �s �  �CYY�M�3�������]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]�f�M��  V��f#�^f;�uj���  f;�u�E�� u9Utj��3�]Ë�U���E������������Dz3��   �E3ɩ�  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������&Q���EQQ�$������U�����  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��f#E�f����E�m�E��Ë�U��QQ�M��t
�-x��]���t����-x��]�������t
�-���]����t	�������؛�� t���]����jh����N��3�9 �tV�E@tH9��t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�� �e��U�E�������e��U�N����A@t�y t$�Ix��������QP�'P��YY���u	��Ë�U��Q�C@V����E�t�{ u�E�>�' �} ~0�E� �M�������E�>�u�?*u�˰?�~����} Ճ? u�E��^�Ë�U���  ���3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������)�����:����������u+��:���    �q:�������� t
�������`p�����7  �F@u^V��L��Y������t���t�ȃ�������� �����A$u����t���t�ȃ������ �����@$��q���3�;��g��������������������������������
  C3�������9������y
  �B�<Xw����0����3����P�j��Y������;�� 
  �$�����������������������������������������������	  �� tJ��t6��t%HHt����	  �������	  �������	  �������	  �������   �	  �������	  ��*u,����������������;��l	  �������������Z	  ������k�
�ʍDЉ������?	  �������4	  ��*u&����������������;��	  ��������		  ������k�
�ʍDЉ�������  ��ItU��htD��lt��w��  ������   ��  �;luC������   �������  �������  ������ �  �<6u�{4u�������� �  �������p  <3u�{2u������������������N  <d�F  <i�>  <o�6  <u�.  <x�&  <X�  ������!�����������P��P�$���Y��������Yt"�����������������C������������������������������  ��d��  �X  ��S��   tL��AtHHt$HHtHH��  �� ǅ����   �������V  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ��u���������������ǅ����   ��  ��X�"  HHt+���  HH��  ��������������  ������t0�G�Ph   ������P������P�7  ����tǅ����   ��G�������ǅ����   �������������|  �����������t;�H��t4������   � ������t�+���ǅ����   �7  !������,  ���������P���Y�  ��p�=  �%  ��e�  ��g��   ��it|��nt.��o��  �������������ǅ����   tl������   �`�������������p��5  ���b��������� tf������f���������ǅ����   �>  ������������@ǅ����
   �������� �  ��  ��W���  ������������@�������   ������������9�����}ǅ����   �ju��gucǅ����   �W9�����~�������������   ~=��������]  V�a��������Y��������t���������������
ǅ�����   ��5<`���������G�������������P��������������������P������������SP�5x����Ћ���������   t������ u������PS�5������YY������gu��u������PS�5������YY�;-u������   C������S�����ǅ����   �������*��s�n���HH�X�������  ������ǅ����'   �������ǅ����   �2���������Qƅ����0������ǅ����   ������   �������� t��������@t�G���G����G���@t��3҉�������@t��|��s����ځ�����   ������ �  ����u3�9�����}ǅ����   ���������   9�����~���������u!������u����������������t-�������RPWS�M�����0�������؋���9~������N뽍E�+�F������   ������������tb��t�΀90tW�������������0@�?If90t����u�+��������(��u����������������I�8 t@��u�+����������������� ��  ��������@t5��   t	ƅ����-���t	ƅ����+���tƅ���� ǅ����   ������+�����+�������������u%���������������� O�0����������t���������������������������P�������2���������YYt.������u%��������������˰0O������������t��ヽ���� ������tu��~q�������������������Pj�E�P������P���1  ����u69�����t.�������������������E�P���������������� YYu��#��������������P�������������]���YY������ |2������t)�������������������� O������������t��߃����� t���������������� Y���������������t���������������r��������� t
�������`p��������M�_^3�[�����Ð98h�c���S��QQ�����U�k�l$���   ���3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|����6�������uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�������h��  ��x����e����>YYt�=`� uV贤��Y��u�6����Y�M�_3�^�S�����]��[Ë�U��UV�uW��H�F��w�� �
�y�B��w�� ��t;�t�_+�^]Ë�U���S�u�M�������]��u#�-���    �L-��8]�t�E��`p������V�u��u$�~-���    �!-���}� t�E��`p������R�E��x uVS�M���YY�1+�W�3�M�QP���������M�QP�������F��t;�t�+���_�}� t�M��ap�^[�Ë�U��3�9,�u'9Eu��,���    �,������]�9Et�]�����P�u�u�������]Ë�U����} SVW��   �u�M�������]��u'�,���    �9,���}� t�E��`p������   �u��tҿ���9}v!�^,���    �,���}� t�E��`p����]�E��x u�uVS�-  ���}� tA�M��ap��8+��3�M�QP��������M�QP������F�Mt��t;�t�+����3�_^[�Ë�U��3�9,�u09Eu��+���    �j+������]�9Et�}���w�]�-  P�u�u�u�������]Ë�U��SV��3�;�u�y+��j^�0�+�����   W9]w�]+��j^�0�+�����u3�9]���A9Mw	�:+��j"�ۋM�����"wɋ�9]t3�C�-�N�؋�3��u��	v��W���0�AC��t;]r�;]r� �� I���I�G;�r�3�_^[]� ��U��}
�Eu
��yjj
�j �u�u�M����]Ë�U���0S3��E�V���]܈]��]��E�   �]�t	�]��E��
�E�   �]��E�P�.  Y����  � �  �Eu�E @ u9E�t�M���E��+ù   ��   �tCHt(Ht �5*������*��j^�0�)������   �M���Et	�E   u��E�   @��U�EjY+�t7+�t*+�t+�t��@u�9U����E���E�   ��E�   ��E�   ��]�E�   #¹   W�   ;�3t(;�t$;�t=   tT=   u-�E�   �T�E�   �K�E�   �B=   t4=   t$;�t)�S)������6)��j^�0��(����_^[���E�   ��E�   �E�E��   ��t�����#M��x�E�   �@t�M�   �M�   �M��   t	}� t	�M�   ��t�M�   ��������;�u!�(���  ��(���    �(��� �`����E�=4aj �u��    �u�E�P�u��u��u�׉E�;�up�M��   �#�;�u+�Et%�e����j �u��E��u�P�u��u��u�׉E�;�u7�6������ ������D0� ��@`P�#(��Y��'��� �E��e  �u���`��uD�6������ ������D0� ��@`��V��'��Y�u�� `��u��'���    렃�u�M�@�	��u�M��u��6�<�����Ѓ����� �Y��Y�M����L��Ѓ����� ����D$� ��M��e�H�M�u~�����  �EtojS�6�p�������;�u�#'���8�   tO�6��]�������j�E�P�6�E� ��������u�}�u�ǙRP�6�(  ��;�t�j j �6������;�t��E���(  � @ � @  �}u�E�#�u	M�	E�E#�;�tD=   t)= @ t"=   t)= @ t"=   t= @ u�E���M�  #�;�u
�E���E� �E   ��  3��E�@�}���  �E��   �#�=   @��   =   �tq;��y  �E�;��n  ��v��v+���[  �E�3�H�  H�G  �E���  j�  jWW�6�8[�����t�WWW�6�'[��#�;������j�E�P�6�!�����;��w�����tj����   �}�﻿ uX�E���   �E�;���   ���i������W���jWW�6�Z������J���WWW�6�Z����#�;���   �����E�%��  =��  u�6��[��Y��$��j^�0�u��_  =��  uWj�6�(�����;�������E��>WW�6��������E�﻿ j[��+�P�D=�P�6��F�������������;�݃��������� ������D$�2M���0������� ������D$�M�������
ʀ}� �u!�Et��ȃ����� ����D� �M��   �#�;�u~�Etx�u�� `j �u��E�jP�u�E�%���P�u�4a;�u4�@`P��#����ȃ����� ����D� ��6�����Y�����6������ �������E��V���SSSSS��"���jh����5��3��}�3��u;���;�u�Q#��j^�0��"�����Y��3�9}��;�t�9}t�E%������@tʉ}��u�u�u�u�E�P���]������E��E������   �E�;�t���5���3��u9}�t(9}�t����������� ��D� ��6����YË�U��j�u�u�u�u�u�!�����]Ë�U���S�u�M������3�9]u8]�t�E��`p�3��  �E�9Xu&�u�u�u�m�����8]���  �M��ap��  9]u&�+"���    ��!��8]�t�E��`p������f  W�};�u&��!���    �!��8]�t�E��`p������7  V�M�	�M�E���D�M�te9]u��D�]���   f����   �U�:�u�]��T����f��E��f��M�f;prf;pwfp�1f;pr+f;pw%fp��U���At	��  ��ʉM�f�u����G�D�M�tG9]u�]��X��M:�t�����f���G�M�f;Hrf;HwfH�1f;Hr+f;Hw%fH��U���At	��  ��ʉM�f�M�f;�u!f;�t	9]�����8]�t�E��`p�3�^_[�����H8]�t��M��ap����U��j �u�u�u�������]Ë�U����} u3���W�u�M������}� u'�u�u�u�Z������}� ��   �M��ap��   S�]��u#� ���    ���8]�t�E��`p������_V�u��u$�����    ����}� t�E��`p������2��M��C�D8t=�} u �3��D8tY�}� t�E��`p�3�^[_�Ê��u3������f���C���F�D:t �} u3����M��t�����f���Ff;�uf��t��} �p�������H�}� t��M��ap�닋�U��j �u�u�u������]Ë�U���8���3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=��O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�����+��;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5��N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3�����A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  ���;����   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�����3�@�   ���e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+����M���Ɂ�   �ً��]���@u�M̋U�Y��
�� u�M̉�M�_3�[�����Ë�U���8���3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=��O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�����+��;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5��N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3�����A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  ���;����   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�����3�@�   ���e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+����M���Ɂ�   �ً��]���@u�M̋U�Y��
�� u�M̉�M�_3�[�����Ë�U���|���3ŉE��E3�V3��E��EFW�E��}��M��u��M��M��M��M��M��M��M�9M$u����    ����3��<  �U�U��< t<	t<
t<uB��S�0�B���  �$�A<�Hπ�wjYJ�ߋM$�	���   �	:ujY������+tHHt���|  ���jY�E� �  뤃e� jY뛍Hωu���v��M$�	���   �	:uj�<+t"<-t:�t�<C�/  <E~
,d<�!  j�Jj넍Hπ��_����M$�	���   �	:�a���:��s����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�h���<+t�<-t��k����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Hπ�wj	��������+t HHt���=���j�����M��jY�Q���j�~����u���B:�t�,1<v�J�&�Hπ�v�:�뿃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�]����B:�}��Q����M��E�O�? t�E�P�u��E�P��  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �!  =�����-  �����`�E�;���  }�ع0��E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k��� �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��   f;��  ���  f;��	  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� ����E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��yB��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  f9E�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �=����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W[�M�_3�^�����ÍI %6w6�6�687p7�7�7�7E8:8�7��U���t���3ŉE��E�U� �  #�S�]�E��A�V#�f�}� W�]��E������E������E����?�E�   t�C-��C �u�}f��u7����   ����   3�f9M�f�����$ �Cf�C0�C 3�@�  f;���   �M3�@f��   �;�u�} t��   @uhĢ�S3�PPPPP���3�f9U�t��   �u9Uu-h���;�u"9Uuh���CjP�h�������u��C�h���CjP�K�������u��C3��k  �ʋ�i�M  �������Ck�M��������3�f�M��ع����`�ۉE�f�U�u�}�M���  ��y�0���`�ۉE�����  �E�T�������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E����E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��yB��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��}����M�����?  ��  f;���  �]��E�3҉U��U��U�U��U�3�#�#Ё� �  �4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��Z���3�3�f9u���H%   � ���E��a���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~K�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m����M��}� ����E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��yB��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t0����)3�f�� �  f9E�f�B0����$ �B�B �s�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�y2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K����C���<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[� ����À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}�f�]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   �é   t��   �}�M����#�#���E;���   ���������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95 ���  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E������Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��3�PPjPjh   @h̢�`���á�����t���tP� `á����3�9������Ë�U���SV�u3�W�};�u;�v�E;�t�3��{�E;�t�������v�����j^�0�p������V�u�M�������E�9X��   f�E��   f;�v6;�t;�vWSV����������� *   �v���� 8]�t�M��ap�_^[��;�t&;�w �V���j"^�0�����8]�t��E��`p��y�����E;�t�    8]��<����E��`p��0����MQSWVj�MQS�]�p�``;�t9]�j����M;�t����@`��z�P���;��s���;��k���WSV�������[�����U��j �u�u�u�u������]����������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U���SVW3�jSS�u�]��]��3���E�#��U���tYjSS�u�w3����#ʃ����tA�u�}+����   ;���   �   Sj�8aP�\`�E���u�����    ����� _^[��h �  �u�  YY�E���|
;�r�����P�u��u��������t6�+��xӅ�uϋu��u��u��   YY�u�j �8aP�D`3��   �=����8u� ����    ����u��;�q|;�skS�u�u�u�|2��#�����D����u設��YP�`�����H��E�#U���u)������    ��������@`��u�#u��������S�u��u��u�2��#���������3��������U��S�]V�u������ ��
����ΊA$�W�y����   ���� @  tP�� �  tB��   t&��   t��   u=�I��
�L1$��⁀���'�I��
�L1$��₀���a��I��
�L1$�!���_^[u� �  ]����% �   @  ]Ë�U��E��u�����    �P���jX]Ë���3�]Ë�U����ES3�VW�E�N@  ��X�X9]�E  3ɉ]���}襥��э<	���ʋU�e ��ى}����֋u����ϋ��M���U�����։0�x�H;�r;U�s�E   �} �t'�u��e �~;�r��s�E   �} �xtA�H�u�e �7;�r;�s�E   �} �XtA�HM��e� ��ɋ��������މH�M�M�M��X�1�2�u�;�r;�s�E�   �}� �t$�S3�;�r��s3�F�ډP��t
�U�B�U�P�M�U�E�} �X�P�����3�9Xu*�P��E���  ��������������P�;�t܉x�x�� �  u0�H��E���  �����������ʉ�H�x�� �  t�f�M�_^f�H
[����%L`�����̋T$�B�J�3��٨�����鲻������̋T$�B�J�3�蹨���`�钻������̋T$�B�J�3�虨������r�������̋T$�B�J�3��y������R�������̋T$�B��t���3��V����h��/����̋T$�B�J�3��9��������������̋T$�B�J�3���������������̋T$�B�� ���3�������p��Ϻ���̋T$�B�J�3��٧���ȵ鲺������̋T$�B�J�3�蹧��� �钺������̋T$�B�J�3�虧���x��r�������̋T$�B�J�3��y����ж�R�������̋T$�B�J�3��Y����(��2�������̋T$�B�J�3��9��������������̋T$�B�J�3������ط��������̋T$�B�J�3�������0��ҹ���M��5����T$�B�J�3��֦���\�鯹���M���P���M����/����T$�B�J�3�訦�����遹���T$�B�J�3�荦���0��f������������hPS�T���YùX��0���h�S�>���Y�h�S�2���Y�h�S�&���Y�h�S����Y�h�S����Y�h�S����Yù��ޘ��h�S�����Y�h�S�����YÃ=�� uK�����t����Q<P�B�Ѓ����    �����tV���`��V��������    ^ùX�阘���|��O�������������r�����r�����rù��Y����	��*���        @� N� ^� n� �� �� �� �� �� ��  � � 4� L� d� t� �� �� �� �� �� �� �� ��  � � &� <� H� R� ^� p� |� �� �� �� �� �� �� �� � &� :� N� j� x� �� �� �� �� �� �� �� 
� � ,� @� L� ^� t� �� �� �� �� �� �� � *� 6� H� V� l� ~� �� �� �� �� ��  �     ��         �R.SDS�R�R�R
SS"S        ��?<LH�        �I�                        ���Q       ~   �� ��     �������N���������������C-DT�!	@-DT�!�?��# � � �p 0�� � ��3D-COAT d:\program files\maxon\cinema 4d r14\plugins\applink_3dcoat\source\applinkdialog.cpp    Start import!   To import a new object? File exists!    export.txt  Folder ..\MyDocuments\3D-CoatV3\Exchange not found! 3D-CoatV3   Exchange    preference.ini  3D-Coat.exe is run! 3D-Coat.exe not found!  open    Start export!       �������N���������������C-DT�!	@-DT�!�?        d:\program files\maxon\cinema 4d r14\plugins\applink_3dcoat\source\applinkexporter.cpp  
       d:\program files\maxon\cinema 4d r14\resource\_api\ge_dynamicarray.h    ]   autopo  curv    prim    alpha   vox retopo  ref uv  ptex    mv  ppp [   # end   v       # begin      vertices
            �?vt   texture vertices
  /   f   usemtl   faces
 g   mtllib  mtl map_    illum 2
    Tr 0.000000
    Ns 50.000000
   Ks  Kd  Ka 0.300000 0.300000 0.300000
  newmtl  No selected objects!    Object "    " has no UVW tag.
UV coordinates can't be exported. Material not found on   object. Default Name    Export object   #Cinema4D Version:  %d.%m.%Y  %H:%M:%S  #File created:  #Wavefront OBJ Export for 3D-Coat
  File     write success! [SkipExport]
   [SkipImport]
         �import.txt  output.obj  obj     �������N���������������C-DT�!	@-DT�!�?�� ���0��T����������string too long invalid string position vector<T> too long  ���P0���� �0��@�0��ios_base::eofbit set    ios_base::failbit set   ios_base::badbit set              Y@��0`p���� 	P	 
�
 ���ܨ``p�P�� 	P	 
����(���� �� �� 00Ppbad locale name Selection   Error on inserting phongTag. Object:    Poly count:     V count:    Create objects...   Memory allocation error for material.   x��"Щ`= 0�6��@�1P	 
 9�9�@�(bad cast        X   ��D    h    can not removed!   normalmap   displacement %f displacement    map_Ks %s   map_Ks  map_Kd %s   map_Kd  Ke %lf %lf %lf  Ke  Ks %lf %lf %lf  Ks  Ka %lf %lf %lf  Ka  Kd %lf %lf %lf  Kd  illum %d    illum   d %lf   d   Ns %lf  Ns  newmtl %s   Open file   .    not found! d:\program files\maxon\cinema 4d r14\plugins\applink_3dcoat\source\applinkimporter.cpp  Nb faces:   Nb Grp:     Wrong face in OBJ file! f   vt  Gathering of data...    �dy���=vt %lf %lf %lf  vt %lf %lf  v %lf %lf %lf   g %s    mtllib %s   Parse file...   Open file:  textures.txt        �������N���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?�pL�K �0�С@�� ��icon_coat.tif   d:\program files\maxon\cinema 4d r14\plugins\applink_3dcoat\source\applinkpreferences.cpp   0��������L          �?x�0U Z�Z�X`U�U�\�������N���������������C-DT�!	@-DT�!�?d:\program files\maxon\cinema 4d r14\resource\_api\c4d_file.cpp �������N���������������C-DT�!	@-DT�!�?     �f@-DT�!	@īP���� �0�@� ����������������     @�@ثP���� �0�@� ���$��� �0�����@�����������d:\program files\maxon\cinema 4d r14\resource\_api\c4d_gui.cpp  l�P���� �0�@� �����P���� �0�@� � �`�p�������������� ��� �Progress Thread 0%  ~   %       �������N���������������C-DT�!	@-DT�!�?d:\program files\maxon\cinema 4d r14\resource\_api\c4d_general.h    %s         �������N���������������C-DT�!	@-DT�!�?�������N���������������C-DT�!	@-DT�!�?����MbP?��� f    d:\program files\maxon\cinema 4d r14\resource\_api\c4d_baseobject.cpp   d:\program files\maxon\cinema 4d r14\resource\_api\c4d_resource.cpp #   M_EDITOR    P���    �������N���������������C-DT�!	@-DT�!�?res     �������N���������������C-DT�!	@-DT�!�?d:\program files\maxon\cinema 4d r14\resource\_api\c4d_pmain.cpp        d:\program files\maxon\cinema 4d r14\resource\_api\c4d_basetime.cpp      �Ngm��C   ����A  4&�k�  4&�kCd������    d:\program files\maxon\cinema 4d r14\resource\_api\c4d_libs\lib_ngon.cpp        �������N���������������C-DT�!	@-DT�!�?d:\program files\maxon\cinema 4d r14\resource\_api\c4d_misc\datastructures\basearray.h  d:\program files\maxon\cinema 4d r14\resource\_api\c4d_basebitmap.cpp   *   ��[�C   ������,�a�@�generic @�������,�a�@�iostream    ��������,�a�@�system  خ������,�a�@�iostream stream error       ��������(�h���t�h���įh����s�s�s�s�s�s�s�s tttttt    r   w   a   rb  wb  ab  r+  w+  a+  r+b w+b a+b          
   !   "   2   *            #   3   +       ���:�\�����Unknown exception   p�����csm�               �                  �?      �?3      3            �      0C       �       ��              fmod         dV��V���V��V�����V�V��V�                                                                                                                                                                                                                                                                                  ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������LC_TIME LC_NUMERIC  LC_MONETARY LC_CTYPE    LC_COLLATE  LC_ALL  �}    ���}����x}��"l}��2�`}��D�X}��^�	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ _., _   ;   =   =;      Visual C++ CRT: Not enough memory to complete call to strerror. H H : m m : s s     d d d d ,   M M M M   d d ,   y y y y   M M / d d / y y     P M     A M     D e c e m b e r     N o v e m b e r     O c t o b e r   S e p t e m b e r   A u g u s t     J u l y     J u n e     A p r i l   M a r c h   F e b r u a r y     J a n u a r y   D e c   N o v   O c t   S e p   A u g   J u l   J u n   M a y   A p r   M a r   F e b   J a n   S a t u r d a y     F r i d a y     T h u r s d a y     W e d n e s d a y   T u e s d a y   M o n d a y     S u n d a y     S a t   F r i   T h u   W e d   T u e   M o n   S u n   HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun K E R N E L 3 2 . D L L     FlsFree FlsSetValue FlsGetValue FlsAlloc    h���e+000   CorExitProcess  m s c o r e e . d l l   p��n��bad exception   r u n t i m e   e r r o r        
     T L O S S   e r r o r  
   S I N G   e r r o r  
     D O M A I N   e r r o r  
     R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
            Ȋ   p�	   �
   Љ   x�   �   Ј   x�   �   ��   H�   ؆   ��   H�   ��    �!   (�x   �y   �z   Ђ�   Ȃ�   ��M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y     
 
     . . .   < p r o g r a m   n a m e   u n k n o w n >     R u n t i m e   E r r o r ! 
 
 P r o g r a m :       �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �            �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow         �������             ��      �@      �               ���5�h!����?      �?            �?5�h!���>@�������             ��      �@      �        united-states   united-kingdom  trinidad & tobago   south-korea south-africa    south korea south africa    slovak  puerto-rico pr-china    pr china    nz  new-zealand hong-kong   holland great britain   england czech   china   britain america usa us  uk  swiss   swedish-finland spanish-venezuela   spanish-uruguay spanish-puerto rico spanish-peru    spanish-paraguay    spanish-panama  spanish-nicaragua   spanish-modern  spanish-mexican spanish-honduras    spanish-guatemala   spanish-el salvador spanish-ecuador spanish-dominican republic  spanish-costa rica  spanish-colombia    spanish-chile   spanish-bolivia spanish-argentina   portuguese-brazilian    norwegian-nynorsk   norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg   german-lichtenstein german-austrian french-swiss    french-luxembourg   french-canadian french-belgian  english-usa english-us  english-uk  english-trinidad y tobago   english-south africa    english-nz  english-jamaica english-ire english-caribbean   english-can english-belize  english-aus english-american    dutch-belgian   chinese-traditional chinese-singapore   chinese-simplified  chinese-hongkong    chinese chi chh canadian    belgian australian  american-english    american english    american        ��ENU ��ENU x�ENU l�ENA d�NLB X�ENC T�ZHH P�ZHI H�CHS 4�ZHH  �CHS �ZHI ��CHT �NLB ԒENU ȒENA ��ENL ��ENC ��ENB ��ENI |�ENJ p�ENZ X�ENS <�ENT 0�ENG $�ENU �ENU �FRB ��FRC �FRL ԑFRS đDEA ��DEC ��DEL ��DES |�ENI l�ITS `�NOR L�NOR 8�NON  �PTB �ESS ��ESB �ESL ؐESO ĐESC ��ESD ��ESF ��ESE p�ESG \�ESH L�ESM <�ESN (�ESI �ESA �ESZ �ESR ��ESU ЏESY ��ESV ��SVF ��DES ��ENG ��ENU ��ENU ��USA ��GBR ��CHN x�CZE p�GBR `�GBR X�NLD L�HKG @�NZL <�NZL 0�CHN $�CHN �PRI �SVK  �ZAF �KOR �ZAF ؎KOR ĎTTO ��GBR ��GBR ��USA ��USA 6-OCP ACP Norwegian-Nynorsk   Illegal byte sequence   Directory not empty Function not implemented    No locks available  Filename too long   Resource deadlock avoided   Result too large    Domain error    Broken pipe Too many links  Read-only file system   Invalid seek    No space left on device File too large  Inappropriate I/O control operation Too many open files Too many open files in system   Invalid argument    Is a directory  Not a directory No such device  Improper link   File exists Resource device Unknown error   Bad address Permission denied   Not enough space    Resource temporarily unavailable    No child processes  Bad file descriptor Exec format error   Arg list too long   No such device or address   Input/output error  Interrupted function call   No such process No such file or directory   Operation not permitted No error    ccs UTF-8   UTF-16LE    UNICODE c c s   U T F - 8   U T F - 1 6 L E     U N I C O D E    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   ->* &   +   -   --  ++  ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __eabi  __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(    ����������|�p�h�`�T�H�c@�8�l~4�0�,�(�$� ����r��� ������d o���������nܞ؞ԞО̞ȞĞ��������������������|�d�X�D�$���ĝ����d�@� ���ܜ̜Ȝ��������x�h�L�,��ܛ����l�H�$���̚��c����l�L�0�GetProcessWindowStation GetUserObjectInformationW   GetLastActivePopup  GetActiveWindow MessageBoxW U S E R 3 2 . D L L     _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          1#QNAN  1#INF   1#IND   1#SNAN  C O N O U T $       ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           ���   RSDS�a��(�F�Z�D)�3   D:\Program Files\MAXON\CINEMA 4D R14\plugins\Applink_3DCoat\obj\applink_cinema4DR14_Win32_Release.pdb                ��           ,�8�T�     �       ����    @   ��        ����    @   p�           ��T�                4���           ����Ԥ    4�       ����    @   ��P�        ����    @   �            �Ԥ                l��           ,�8�Ԥ    l�       ����    @   �            ��h�           x���    ��        ����    @   h�           ������    ��       ����    @   ��           ����    ��       ����    @   ԥ            �� �           0�<�X�    ��       ����    @    ��       ����    @   t�           ����    �        ����    @   t�           $���           ̦���T�p�    $�       ����    @   ��`�              P   �           (�8�<�X�    `�       ����    @   ���              @    ��              @   t�            `��            ����           ħԧ���    ��       ����    @   ��            ���           �$�8�Ԥ    ��       ����    @   �            ��T�           d�x�$�8�Ԥ    ��       ����    @   T�            ����           ����    ��        ����    @   ��            8��            ����    8�       ����    @   �            ��<�           L�\�����    ��       ����    @   <�    X       ����           �������T�p�    ��       ����    @   ��            ���           �� ���    ��       ����    @   �    h       T�0�           @�X����T�p�    T�       ����    @   0�           ������    ��       ����    @   t���        ����    @   Ȫ           ت��                ����           ������    ��       ����    @   ��            ��D�           T�\�    ��        ����    @   D�            ���           ����\�    �       ����    @   ��            �p�            0��           ���T�    0�       ����    @   �            L�8�           H�P�    L�        ����    @   8�            h���           ����T�    h�       ����    @   ��            ��̬           ܬ���T�    ��       ����    @   ̬            ���           ,�4�    ��        ����    @   �            ��Ȫ            ��x�           ����    ��        ����    @   x�            ����           Эܭ��    ��       ����    @   ��            ���           �$�    ��        ����    @   �            �T�           d�p�$�    �       ����    @   T�            D���           ����$�    D�       ����    @   ��            p��           ���p�$�    p�       ����    @   �            ��<�           L�X�Ԥ    ��       ����    @   <�            ����           ����X�Ԥ    ��       ����    @   ��            ��د           ���X�Ԥ    ��       ����    @   د            ��(�           8�@�    ��        ����    @   (�            P��            8���           ����Ԥ    8�       ����    @   ��            ��а           ��Ԥ    ��       ����    @   а        c m �\ �� �� `P �P �P �P �P  Q  Q @Q `Q �Q �Q �Q �Q  R  R @R cR �R �R                     P�     ��   ����    4�    ����       @    P�    ����       ��    P    �   ���0���    ��    ����       `    ��    ����       `    l�    ����       @    P    \�   0���            y            ����    ����                  "�   ��   ̲                            x�              h�    ��    �   ���    8�    ����       ��            �!����    ����                  ,�"�   <�   L�                            �$����    ����                  ��"�   ��   ��                            �%����    ����                  ܳ"�   �   ��                            �'����    ����                  4�"�   D�   T�                            O(����    ����                  ��"�   ��   ��                            �+����    ����                  �"�   ��   �                            �.����    ����                  <�"�   L�   \�                            �0����    ����                  ��"�   ��   ��                            �<����    ����                  �"�   ��   �                            4?����    ����                  D�"�   T�   d�                            �C����    ����                  ��"�   ��   ��                            �F����    ����                  ��"�   �   �                            �T����    ����                  L�"�   \�   l�                            W����    ����                  ��"�   ��   ķ                            8X����    ����                  ��"�   �   �                ����[R"�   T�                       ����~R    �R"�   ��                           ��    ����       ��    ��    �   �����    ��    ����       ��    ��    �   ,�����    ��    ����       K�����    ����    ����    �    ����    ����    ����    �    ����    ����    ����        ����    ����    ����    E
        
����    ����    ����    �
    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    6    ����    ����    ����    Q    ����    ����    ����    �    ����    ����    ����Sd    ����    ����    ����    (    ����    ����    ����    �3        �3        �3    ����    ����    ����    �5    ����    ����    ����    �6    ����    ����    ����    u8    ����    ����    ����    �;    ����    ����    ����    �?    ����    ����    ����    C    ����    ����    ����    DD����    SD����    ����    ����    F����    F����    ����    ����    �`    ����    ����    ����    &c    ����    ����    ����    �d    ����    ����    ����    �l    ����    ����    ����    �m    ����    ����    ����    �o    dono����    ����    ����JpSp@           ,q����    ����                  ��"�   �   �                   ����    ����    ����    dr    �q�q����    ����    ����KtOt    ����    ����    �����t�t    n    ̽   ؽ��    ��    ����       �y    ����    ����    �����z{    ����    ����    ����N{R{    ����    ����    ����    y    ����    ����    ����    �    ����    ����    ����    G�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    9�    ����    ����    ����k�~�    ����    ����    ����    ��    ����    ����    ����    ��        ������    ����    ������    ����    ����    ����    '��         ��  ` 8�         �� @a                     @� N� ^� n� �� �� �� �� �� ��  � � 4� L� d� t� �� �� �� �� �� �� �� ��  � � &� <� H� R� ^� p� |� �� �� �� �� �� �� �� � &� :� N� j� x� �� �� �� �� �� �� �� 
� � ,� @� L� ^� t� �� �� �� �� �� �� � *� 6� H� V� l� ~� �� �� �� �� ��  �     ��     R CloseHandle �Process32Next ZModule32First �Process32First  � CreateToolhelp32Snapshot  KERNEL32.dll   ShellExecuteExA SHELL32.dll �InterlockedIncrement  �InterlockedDecrement  �Sleep �InitializeCriticalSection � DeleteCriticalSection � EnterCriticalSection  9LeaveCriticalSection  � EncodePointer � DecodePointer GetLastError  �HeapFree  �RaiseException  RtlUnwind � DeleteFileA �GetCurrentThreadId  �GetCommandLineA �HeapAlloc WideCharToMultiByte -LCMapStringW  gMultiByteToWideChar rGetCPInfo hGetACP  7GetOEMCP  
IsValidCodePage �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree GetModuleHandleW  sSetLastError  EGetProcAddress  �UnhandledExceptionFilter  �SetUnhandledExceptionFilter  IsDebuggerPresent �TerminateProcess  �GetCurrentProcess IsProcessorFeaturePresent �HeapCreate  �HeapDestroy oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW ExitProcess %WriteFile �GetConsoleCP  �GetConsoleMode  WFlushFileBuffers  �ReadFile  fSetFilePointer  GetModuleFileNameW  GetLocaleInfoW  GetModuleFileNameA  aFreeEnvironmentStringsW �GetEnvironmentStringsW  �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime �HeapSize  iGetStringTypeW  �HeapReAlloc �GetUserDefaultLCID  GetLocaleInfoA  EnumSystemLocalesA  IsValidLocale ?LoadLibraryW  $WriteConsoleW �SetStdHandle  � CreateFileA � CreateFileW SSetEndOfFile  JGetProcessHeap                    ���Q    R�          H� L� P� �� j�   applink_cinema4DR14.cdl c4d_main                                                                                                                                              Xt    .?AVApplinkDialog@@ Xt    .?AVGeDialog@@  Xt    .?AVbad_alloc@std@@ Xt    .?AVexception@std@@ Xt    .?AVruntime_error@std@@ Xt    .?AVfacet@locale@std@@  Xt    .?AVcodecvt_base@std@@  Xt    .?AUctype_base@std@@    Xt    .?AVios_base@std@@  Xt    .?AV?$_Iosb@H@std@@ Xt    .?AV?$basic_istream@DU?$char_traits@D@std@@@std@@   Xt    .?AV?$basic_ios@DU?$char_traits@D@std@@@std@@   Xt    .?AV?$ctype@D@std@@ Xt    .?AVsystem_error@std@@  Xt    .?AVfailure@ios_base@std@@  Xt    .?AV?$basic_streambuf@DU?$char_traits@D@std@@@std@@     Xt    .?AV?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    Xt    .?AV?$codecvt@DDH@std@@ Xt    .?AV?$basic_istringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    Xt    .?AV?$basic_filebuf@DU?$char_traits@D@std@@@std@@   Xt    .?AVbad_cast@std@@  Xt    .?AV?$basic_ifstream@DU?$char_traits@D@std@@@std@@  Xt    .?AVCommandData@@   Xt    .?AVBaseData@@  Xt    .?AVApplinkPreferences@@    Xt    .?AVTriangulator@@  Xt    .?AVCTriangulator@TRIANGULATOR@@    Xt    .?AVGeModalDialog@@ Xt    .?AVGeUserArea@@    Xt    .?AVSubDialog@@ Xt    .?AViCustomGui@@    Xt    .?AVNeighbor@@  Xt    .?AVC4DThread@@ ����Xt    .?AV_Locimp@locale@std@@    Xt    .?AVerror_category@std@@    Xt    .?AV_Generic_error_category@std@@   Xt    .?AV_Iostream_error_category@std@@  Xt    .?AV_System_error_category@std@@     s�r(ssLs�r@s   Xt    .?AVlogic_error@std@@   Xt    .?AVlength_error@std@@  Xt    .?AVout_of_range@std@@      
       Copyright (c) 1992-2004 by P.J. Plauger, licensed by Dinkumware, Ltd. ALL RIGHTS RESERVED.              Xt    .?AVtype_info@@ N�@���Du�  s�          @�    @�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             sqrt    PvRxTx                                                                                                                                                                                                                                                                                                                                                               abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     p��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����C   � ����������܁ԁȁ��������������������������|�x�p�d�\�T���L�D�<�0�(��������܀	         Ԁ̀Ā������������t�`�L�<�(� ���� ������������ ��tdP@,�~�~�~                                                                                           ��            ��            ��            ��            ��                              8�        Pv�zX|�� � �p���������                                     	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 /�/�/�/�/�/�/�/�/�/������
                                                                                                                                                                                                                                                                                                                                                    Xt    .?AVbad_exception@std@@ ?                 .          .   .   0�d�d�d�d�d�d�d�d�d�4�h�h�h�h�h�h�h�8�    ̙������l�X�<�(�� ��Ș��������t�h�X�H�8�(����������������l�\�P�@�,���������̖������+                                                                                                                                                                                                                        �            �&         ��   �   �   �   0�   (�!    �   ܍   ԍ   č   �   �   ��   ��    ��   ��   ��   �   ��    �   ��   �   �   �"   ܡ#   ء$   ԡ%   ̡&   ��      �      ���������              �       �D        � 0     H�8�   ���5      @   �  �   ����             ����         �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                                                                                                                                                                                                                                                                                       �   40E0t0�0�0�0�01J142]233A3S3f3�3�3�3�3	44,4J4\4n4�4�4�4�4�4�4�6�7�7�7�7�78Q8^8�8�8�899+9<9N9_9h9�9�9�9�9�9�9�9
::1:E:X:j:{:�:�:�:;`;�;�;�;�;<4<h<�<�<�<=I=�=�=�=>P>b>t>?�?�?�?�?�?      �   �0�0�0�011*1M1a1s1�1�1�1�1�1�12<2O2W2n2�2�2�2�23&373I3]3�35535C5�5�5�5�56�6�6�6�6�6�67	7y7�7�78B8Y8y8�89F9�9�9:5:J:R:i:�:�:�:�:;;,;:;�;<<+<D<K<d<|<�<�<�<�<	=+=D=\=u=�=�=�=�=�=>8>J>\>n>v>�>�>�>�>�>�>�>�>�>�>�>�>�> 0  T  
2$262?2P2b2k2�2�2�2�2�2�2�23!363J3c3u3�3�3�3�3�3	44$464H4P4e4z4�4�4�4�4�4�45)5T5i55�5�5�5�5 66+6?6[6m6�6�6�6�6�6�6	7767M7i7~7�7�7�7�7�78&8<8M8b8w8�8�8�8�8�8�8�89%9:9R9�9�9�9�9�9�9�9 ::&:;:O:e:y:�:�:�:�:�:�:;";4;E;Z;r;�;�;�;�;�;<"<1<D<W<j<|<�<�<�<�<�<�<='=9=K=\=q=�=�=�=�=�=�=>>->B>J>_>w>�>�>�>�>?)?@?Y?s?�?�?�?�?�?   @  d  0&0E0Z0u0�0�0�0�0�01&1A1X1w1�1�1�1�1�12272M2^2s2�2�2�2�2�2�233-3B3Z3u3�3�3�3�3�3�3�34$4,4A4Y4s4�4�4�4�4
5"5;5R5�5�5�5�5�5�5	6(6=6X6o6�6�6�6�6�6	7$7;7Z7o7�7�7�7�7�78&8?8S8h8}8�8�8�8�8�8�89"979O9g9�9�9�9�9�9�9�9�9::3:H:T:�:�:�:�:�:;,;D;n;�;�;�;�;�;�;<(<C<Z<y<�<�<�<�<�<=&=E=Z=u=�=�=�=�=�=>*>>>S>h>|>�>�>�>�>�>�>?"?:?R??�?�?�?�?�?�?�? P  l  0
0070C0y0�0�0�0�01141Z1q1�1�1�1�1�1�12212M2_2t2�2�2�2�2�23343K3j33�3�3�3�3�34$454G4Y4m4�4�4�4�4�4�4�455J5_5h5y5�5�5�5�5�5�5�56&6?6Q6f6z6�6�6�6�6�6�67"7G7z7�7�7�7;8M8_8y8�8�8�8�8�8�8&999K9_99�9�9�9�9:::/:A:J:b:t:�:�:�:�:�:�:	;;0;B;T;e;|;�;�;�;�;<!<*<@<U<k<}<�<�<�<�<�<�<=+=A=R=d=v=�=�=�=�=�=>>$>9>�>�>�>�>�>�>�>?'?0?B?[?o?�?�?�?�?�?�? `  l  00-0?0Z0y0�0�0�0�0�01&1;1D1X1t1�1�1�1�1�12 2L2^2p2x2�2�2�2�2�2
3323N3�3�3�3�3�3�3�34@4R4d4m4�4�4�4�4�4�4�45535L5^5s5�5�5�5�5�5�5�56)6N6b6w6�6�6�6�6�67707Z7l7~7�7�7�7�7�7�7�78(8=8X8~8�8�8�8�899+9=9U9i9�9�9�9�9�9�9	: :<:N:f:z:�:�:�:�:�:�:;&;8;L;^;p;�;�;�;�;�;�;�;�<�<�<�<�<�<�< ==*=C=U=j=~=�=�=�=�=�=�=>>6>H>[>o>�>�>�>�>�>�>?9?J?�?�?�?�?�? p  $  0/0a0r0�0�0�081M1b1w11�1�1�1�1�1�12202F2Z2v2�2�2�2�2�2�23%3:3C3[3s3�3�3�3�34%444Z4o4�4�4�4�4�4�455535L5`5|5�5�5�5�5�5�56�6�6�6�67L7]7�7�7�7�7�78(8:8M8�8�8�8�8�8909C9�9�9�9�9:?:h:�:�:>;�;�;�;�;�;<<0<i<{<�<�<�<�<�<= =H=Z==�=�=�=�=�=>>'>j>{>�>�>�>?2?C?U?g?p?�?�?�?   �  �   	00+040F0W0s0�0�0�0�0�0�0
1!1>1P1b1j1|1�1�1�1�1�122*2>2U2}2�2�2�2
3343<3k3�3�3�3�3�344>4�45Q5o5�56A6Y6�6�6�6�6�6�67u7�7�78 8?8^8B9�=�=�>   �  �   31f1�1�1�12J2^2s2�2�2�2�2"3H3Y3l3u3�3�3�3�3�3�3�34434G4j4|4�4�4�4�45505B5b5R6`6!767�7�7R8`899�9�9�9:p:~:8;=;�<�<
=p>~>#?-?I? �  �   �0�0�0t1�1�1�1R2R3�45#5=5U5n5�5�5�5�56O6�6�6�67 7,7W7t7�7878W8�8�8�8949N9`9l9�9�9:S:�:�:�:;.;@;L;w;�;�;3<e<�<�<�<!=T=n=�=�=�=�='>s>�>�>?M?z?�?   �  �   0+0?0T0�0�0 1P1q1�1�1�1�1�1�12222G2[2w2�2�2�2�2�23"3*3C3Y3o3�3�3�3�3�34#484Q4�6�67 757=7S7j7�7�7�7�7�78#8S8q8�8�89<9Q9Y9u9�9�9�9�9�9 ::;:O:d:y:�:;5;_;�;�;E=�=>&>8>e> �  �   0*0V0l0t0�0!161K1S1h1}1�1�1�1�1�12+2B2n2�2�2�2�2�23$383M3V3k3�3�3�3�3�3�3404G4s4�4�4�4�4E5�5�5�5�5�56<6U6w6�6�6�6�67=7Y7�7�7�7�78.8[8y8�8�8U9k9s9�9:4:I:R:f:{:�:�:�:;;.;V;h;�;�;�;�;�;G<\<q<�<�<2=G=g=�=�=>b>v>�>�>?)?[?~?�? �  �   0#0+0@0U0^0r0�0�0�0�0�01&1=1i1~1�1�1�1�1�12r2~2�2�2�35�5�5�5�5�566)6B6V6u6�6�6�6�6�6737G7\7q7�7�7�7�7 8a8�8�8]9s;�;�;�;<,<V<[<�<=%=Z=o=�=%>9>N>a>w>�>�>�>�>�>?7?L?`?�?�?   �  �   /0:0j0(1<1P1Y1n1�1�1�1�1�1�12!262Q2h2�2�2�2�2�23k3�3�3�3�3�3�3�3�3414H4g4|4�4�4�4�455-5A5s5�5�5�5+6M6�6�6"878P8l8�89~9�9�9f:n:x:�:�:�:%;H;{;�;�;�=#>   �  �   b1�2�2�23'3�3�3�3!4�4�4z5�5�5�5�5�5656L6a6v6�6�6�6�6�6
77b7w7�7�7�7�7	88c8w8�8�8�8y9�9�9�9�9�9�9:':>:X:m:�:�:�:�:�:
;;M;y;�;�;�;�;�;�;<#<=<R<n<�<�<�<�<�<=�=�=�=�=�=�=>>:>O>m>�>�>�>�>�>?+???T?i?   x   0Q1a1�1�1�1�1�1	2222G2d2w233A3W3l3�3�3�3�34�5�5�5�5�5�566.6Q6r6r7�7�7�7�:�:(;.;�<�<S=Y=�=�=�=>�>�>?
?h?    T   Q0�0�0�1-2�3�3B4M4�4�455�5�5�6�6�6�6{7�7�7w8�8�8�;�=>�>R?X?m?u?{?�?�?�?�?   d   	0�061F1�1�1�1�1�2�2�2�2�3�3�4&585X5B6H6]6e6k6p6�6�6�6�667H7�7�7�8�8�9�9f:x:�;�<�=F>[>??   0 @    161H1W1i1z1�1�3�3�3D4X4'5�6�9�9�:�:�;�;�;<l=�=F>X>y>   @ H   %1,181�1�1�122Z2�23(3�4�5�5�5�6�:;;';c;�;�;�;�;�;I<�<q>�?   P d   �23Z3r3�3�34484�466�6�6f7x7�7|8�<�<�<�<�<�<=D=d=�=�=>�>�>�>�>??4?E?S?t?�?�?�?�?�?�? ` $  0$0D0d0�0�0�0�0�0�0141L1`1o11�1�1�1�1�1�12C2V2j2z2�2�2�2�2�23$3<3P3`3�3�3�3�344'4D4t4�4�4�45545a5t5�5�5�5�5646T6q6�6�6�6�6�67$7D7d7�7�7�7�78858d8~8�8�8�8�89-9D9�9�9�9�9�9:g:�:�:�:�:�:�:H;�;�;�;�;<D<d<�<�<�<�<=$=D=d=�=�=�=�=>>$>Q>d>>�>�>�>�>�>?? ?A?d?�?�?�?�?�?�? p (  0040O0]0k0z0�0�0�0�0141T1t1�1�1�12 212M2w2�2�2�2�2�2343T3t3�3�3�3�3�34404T4n4�4�4�4�4�4�4555L5]5k5�5�5�5�5�566%656F6�6�6�6�67$7T7a7q7�7�7�7�78$8D8d8�8�8�8�89$9D9d9�9�9�9�9:$:D:d:�:�:�: ;$;D;d;�;�;�;�;<$<D<d<�<�<�<�<=$=D=d=�=�=�=�=>$>D>d>�>�>�>�>�>?$?A?Q?a?t?�?�?�?�?�?   � �   $0D0i0�0�0�01�1�1�142T2n2v2�2�2�2313D3W3x3�3�3�344D4d4�4�4�4�4$565d5�5�5\6�6�6�6�677w7E8J8U8x8�8�8�8�89A9t9�9�91:d:�:�:�:*;V;k;�;�;<K<�<�<�< =P=�=�=�=�=�=>6>M>w>�>�>�>?1?P?l?�?�?�? � �   010k0�0�0�0�01G1q1�1�1�122g2�2�2�2�2*3�3�3�3�3U4�4�4K5�5�5�5(6k6�6�6	7#7l7�7�7868Q8�8�8�89d9�9D:�:�:$;=;a;s;�;�;�;�;=<�<�<=a=�=�=�=2>k>�>�>�>�>�>1?j?�?�? � t   t0�01`1�1�1@2�2�2S3�34S4�45s5�536�6�6S7�78c8�8#9�9�9:�:�:@;p;�;�;<@<p<�<�<=]=�=�=�=�=$>^>�>�>?k?�?   � �   0N0�0�0121T1�1�1242t2�2�2%3E3^3�3�3U4Z4e4{4�4�4�4�4h5�5�536�6F7�7�7�7�7�7�7�7�7�7�7�8�8�8�8�8 99999�9�9�9:/:B:^:�:�:�:�:;$;d;�;�;�;<4<d<�<�<=D=d=�=�=�=>+>H>Z>�>?$?T?�?�?�?�?   � �   $0T0�0�0�0�0�01!131G1d1t1�1�1�1�1�12222O2[2f2�2�2313Q3t3�3�34D4t4�4�45D5t5�5�56D6^6747u7�7�7�7P8�8�8�8�8�9�9H:u:z:�:�:�:�:�:1;�;�;�;�;�;
<4<T<t<�<8=�=>D>t>�>�>?'?E?_?|?   � �   #0S0q0�0�0�0!161J1_1�1�1�112h2m2y2�2�2�234314o4�4�4�4�4�45W5x5�5�5�5�5(6L6e6~6�6�67 7G7�7�7�7�7�7�78.8L8j8�8�8�8,9^9�9�9(:�:�:;4;c;�;�;�;�;B<t<�<�<�<=+===Y=g=�=�=�=�=�=>>'>?>T>o>�>�>�>�>�>�>? � �   �0�1�1$2t2�2I3�34�4�4�4(5I5u5�5	6�6�6�7�7�7�7�7�7	8808B8V8s8�8�8�8999M9i9�9�9�9:!:-:B:U:i:{:�:�:�:�:�:;;9;P;�;�;�;�;�;[=e=�=�=>#>A>a>t>�>�>�>?4?O?o?�?�?�?�? � �   040t0�0�0�0�01D1d1�1�1�1212T2�2�2�2�2343T3t3�3�3�3�3414D4d4�4�4�4.5N5c5�56a6�6�6X7z7�78:8]8�8�89~9�9�93:\:�:�:�:$;�;�;<�<�<�<c=�=�=.>N>c>�>L?w?�?�?   �   Q0w0�0�0Q1�132\2�2�2333�3�3�314G4�455�5�5�5�5646T6k6�6�6�67A7a7�7�7�7�78G8q8�8�8�8979K9j9�9�9�9:4:Q:q:�:.;3;8;=;_;�;�;�;�;<$<D<d<�<�<�<=4=T=q=�=�=�=�=�=2>`>�>�>?0?^?�?�?�?�?  �   040d0�0�0�0�0$1D1t1�1�1�1$2D2d2�2�2�2�23$363Q3d3�3�3�3�3�34$4a4q4�4�4�45$5D5a5t5�5�5�5�5�5646T6t6�6�6�67$7A7T7t7�7�7�7�78d8�8�8�8�8949T9t9�9�9�9�9:W:�:�:;S;�;�;<$<T<�<�<�<�<=!=1=D=d=�=�=�=�=>->f>�>�>�>�>?&?T?t?�?�?�?       00D0b0v0�0�0�0�0141T1�1�1�1�1�1242Z2�2�2�2�2�2�23"3D3^3r3�3�3�3�3�34D4X4�4�4�4�4�4505I5W5f5�5�5�5�56,6@6Y6g6v6�6�6�67$787N7�7�7�7�788.8d8�8�8�8�8949T9t9�9�9�9�9::T:t:�:�:�:�:;4;T;t;�;�;�;�;�;<$<T<q<�<�<�<�<�<�<==/=H=Z=l=�=d>�>�>�>5?r?�?�? 0 �   E0u0�0�01X1�1�12O2�2�23B3u3�34R4�4�45E5u5�5�5%6U6�6�657u7�7�78@8T8d8�8�89U9�9�9%:e:�:;);Q;y;�;�;�;�;<*<U<y<�<�<=?=�=�=�=%>M>v>�>�>?C?h?�?�?�? @ �   0=0x0�0�0!1�1�1�1�12$2D2d2�2�2�2�2�2�23!343T3t3�3�3�3�3414T4q4�4�4�45$5D5d5�5�5�56!616D6d6�6�6�6�6�6!7?7d7�7�7�7�7%8=8L8q8�8�8�8�8�8	99d9�9�9�9:$:Q:t:�:�:�:;T;�;�;4<T<t<�<�<�<�<=4=d=t=�=�=�=>D>d>�>�>�>?1?T?�?�?�? P �   0$0g0�0�0�0�0111Q1q1�1�1�1�1212Q2q2�2�2�2�23A3_3�3�3�3�34$4A4a4�4�4�4�45$5D5a5�5�5�5�5646T6q6�6�6�67�7�78D8d8�8�8�89$9A9d9�9�9�9:4:d:�:�:�:B;a;�;�;�;�;<D<q<�<�<�<�<=D=t=�=�=�=>4>T>�>�>�>�>�>?A?P?t?�?   ` �   40a0t0�0�0�01A1a1�1�1�12!2A2d2�2�2�2$3T3�3�3�34Z4�4�4�4515T5�5�5�5�5�56-6j6�6�67$7J7�7�78 8�89Q9e9z9�9�9�9:S:v:�:�:;$;D;�;�;@<�<�<�<�<=I=s=�=�=�=�=>3>T>�>�>�>�>?4?T?�?�?�? p �   0A0a0�0�0�0�01d1�1�1�12422�2�2�2!3>3h3�3�3�3�34,4L4f4�4�4�4�45"5_5s5�5�5�5606U6o6�6�6w7�7�7�78 8>8�8�:A=Z=�=�=�=�=!>^>y> � �   (0,00040�1�152�34�4�4e5�5�5�5�6�67t7�7�7�788A8t8�8�8�8	9%9F9v9�9�9�9�9:1:A:]:�:�:�:�:�:(;];k;z;�;�;�;G>�>?S?�?�?   � H  0*090d0m0z0�0�0�0�0�0�0�01161U1g1�1�1�1�1�122272I2[2m22�2�2�2�2�23$363H3Q3o3�3�3�3�3�34"4/4G4Y4k4}4�4�4�4�4�45545F5X5a55�5�5�5�5�5�56>6T6p6�6�6�6�6�6�6�677/787V7t7�7�7�7�7�7�788@8V8r8�8�8�8�8�8�89"949=9[9|9�9�9�9�9�9:1:�:�:�:�:�:�:; ;1;:;M;�;�;�;�;
<<.<T<q<�<�<�<==m=�=�=�=�=�=�=">?>v>�>$?9?[?�?�? � �   0!010D0�0�0�0�0�01$1A1T1t1�123	3333%3,333:3h3�3�3�3�3�45�6�6�6K7�7�7�7�7�7�7�788888$8+82898@8�9�9�9�9�9:!:;:o:�:�:�:�:�:�:�:�:�:�:';G;�;<U<l<�<�<�<�<=6=D=�=�=>!>D>a>�>�>�>U?a?k?q?v?�?�?�?�?   � 8   0A0T0q0�0�0�011(13181d1{1�1�1	212Q2q2�2�2�6   � h   �0�01U1�1�1%2e2�2�23E3�3�3�354u4�4�4"5R5�5�5�5%6e6�67E7�7�78U8�89e9�9�95:<7<�>(?,?0?4?8?   � �   0)0H0V0�0�011�1�122W2e2|3�3�3�3 4.4C4Q455A5d5�5�5�5�56&6Q6t6�6�6�6747d7�7�7�7�78D8t8�8�8�8949Q9q9�9�9�9�9$:V:k:�:;$;T;�;�;�;�=�=�= >�>? � �   �0�0�0141T1�1�1�1�1�1�12D2t2�2�2�2�23$3A3d3�3�3�3�3�45j5o5�5�607E7U7�788n899C9�9�9�9T:�:<"<,<<<H<N<X<h<�<�<�<�< =+=<=H=P=V=e=n=�=�=�=�>�>�>??+?Q??�?�?�?�?�?�? � �   �0�0�0�1�1�1�1262A2]2�354A4�4�4�4�4�4	5555%5,52595E5�5q6y6�6�6�6�8L9�9�9�9�9�9�9�9�9�9::::::!:':+:1:5:�:�:�:�:�:�:�:�:;?;];d;h;l;p;t;x;|;�;�;�;�;�;�;B<M<h<o<t<x<|<�<�<�< ========f=l=p=t=x=�==>�>�>�>�>?Z?�?�?�?�?�?�?�?�?     �   0-04080<0@0D0H0L0P0�0�0�0�0�01181?1D1H1L1m1�1�1�1�1�1�1�1�1�1�162<2@2D2H2_3e3w3�3�3�3;4B4d4k4�4/565X5_5�5�5!6�67707?7L7X7h7o7~7�7�7�7�7�7�7�7 8S8b8k8�8�8w9�9�9�9:Q:�:Y;�;�<�<�<-?M?    �   S1�2�3f4p45�5�56W6\6f6�6�6�6�6�60767<7Q7�7�7�7
878�8�8�8�829z9�9:1:::B:b:~:;;$;�;�;�;�;�;�;�;�;Q<[<�<�<==/=C=�=%>�>s?{?�?�?     p   g0s0�0�0j1v1�1�12�2�4p5�5�5�5�5�5�5�56(646k6t6�6�6�6�677 7N7�7|89a9�9�9�9�9�9;:V:g:�:;�;�<6=:?j?�? 0 �   00p0�01O1W1�2333a3k3w3�3�3�3�4�4 5�5f6�67-781868j9�9�9.;?;y;�;�;�;�;�;�;�;�;<<0<T<�<�<�<C=`=�=>7>�>�>�>�>�> ???8?T?]?c?l?q?�?�?�?�?�? @ ,  A0�0�0,1�12�2�2�2�2)303<3B3N3T3]3c3l3x3~3�3�3�3�3�3�3�3�3�3�3"4b4h4�4�4�4�4�4�4l5�5�5�5�5%656;6G6M6]6c6i6x6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6
77777$7)7/747C7Y7_7g7l7t7y7�7�7�7�7�7�7�7�7�7�7-8?89)969t9{9�9�9�9�9
::�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;	;;;";-;9;>;N;S;Y;_;u;|;@<E<�>#?i?   P `   �4�5!7'7-7r8~8�8�8�8N9e9�9�9�9 :e:l:�:�:�:�:;3;W;�;�;�;�;�;<%<J<�<�<�<�=�=�=>^>s?z?�? ` �   0@0I0p0}0�0�0�0�0�0�0�0k1s1�1�1�1�1�1�1�1�1�1�12#2+2;2A2R2�2�2�2�2�2�23�3�3�3�3�3�3�3�3�34*40494L4p4�45$5;5�5=6]6M7v7�7=9:�:;.;o;�;+<]<�<�<)=I==�=>>�> p <   
0�0G1�2b4�7�7�7�7�9�:-;8;>;c;i;n;�;;<=�=?�?�?�?   � (   0G0o0	1F1P1h1�1�1�13�3�3�3�:�: � �   K5R5p5�5�5�5�5�56!6'656i6v6�6�6�6%7S7}7�7�89&9.9=9u99�9�9�9�9�9�;�;�;�;�;�;G<M<i<�<�<�<�<�<=#=�>�>�>�>�>�>?4?<?N?[?a?�?�?�?�?   � �   0L0�0�0�0�0�0�0�011&1Q1l1s1|1�1�1�1�1�1�1�1�1222 2$2(2,2024282<2@2D2L2Q2i2�2 4&4D4�4�4�5�5�5�5�5�5�6@7�7\89:,:=:E:U:f:,;O;�;�<�<�<===Q=i= � D   n9�9�9�9:":4:k:�;�;�;�;�;�;J<\<n<�<�<�<�<�<�<�<�<="=\=�?   � D   B0S0}2�2�2�2�2�2k3�3,4m4�4>6{657>7�7�7�78a8j8�8�8�89&9>   � P   ]>a>e>i>m>q>u>y>}>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>!?'?5?   � t   �01$1C1�1�1�1�1)292c2t2�2�2�2�2�23!3,4�4�4�4�4�4$56�687=7B7G7W7�7�7�7�7�788&8+82878E8�8�8�869�:�:�;�=�? � �   0�1C2M233�3�3i4s45Q5�5�5�6�6�671777�7�7�7	8858�8K9�9�9�9:R:e:}:�:�:;1;M;z;�;�;�;�;�;7<I<�<�<�<�<==W=�=>>�>�>�>�?�?�?�?     h   000 0&00060@0F0P0Y0d0i0r0|0�0�0�0�0�2�23)3?3�3�6+8F8\8r8z8�8�9`:�:�:E;i={=�=�=�=�=�=�>f?�?�?  4   
0040I3?4�56B6c6G8�:�:�:�:�:�:�:�:�:�; =)>   H   �0{1�1�12*2=2O2�2�2�5�5�56%6/6F6k6�6;7�:;s<{<,=>�>�>L?R?`?�? 0 T   0M0�0�1�1}2^3�3�3�4�4�4M5d5�5!6�8�8A<E<I<M<Q<U<Y<]<a<e<i<m<z<<=d=t=�=�=>   @ ,   8�9�9�9�9�9�9�9�:;<<C<�<�<!=N=�=e> P h   V0r0�0�0�0�0121U1r1�1�1�1�1222R2u2�2�2�2�2�2�2�233#3/393E3R3Z3d3v3�3�3�3�3�3�3�3�3�3�3�3�3�3 ` �  L1P1T1X1\1`1d1h1l1x1|1�1�1�1�1�1�1�1 22222222�6�6�6�6�6�6�6�6 777777T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9�9�9<<<< <$<(<,<0<4<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >$>h>l>p>t>x>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�?�?�? p �   �0�0�1�1�1�1�1�2�2�2�2�2�2�2�2�2�2 333333$3(3,3034383<3H3L3P3T3X3\3`3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3T4X4\4`4d4h4�4�4�45555 5$5(5,5054585<5@5D5H5L5�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= � @   P2T2�2�2�2�2,;4;<;D;L;T;\;d;l;t;|;�;�;�;�;�;�;�;�;�;�;�; � �   �3�3�3�3�3�3�3�3�3�3 4444 4(40484@4H4P4X4`4h4p4x4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 5555 5(50585@5H5P5X5`5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 6666 6(60686@6H6P6X6`6h6�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? � �   00000000 0$0(0,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1014181<1@1|3�344(4,40484P4T4l4|4�4�4�4�4�4�4�4�4�4�4�4 555(5,50585P5`5d5t5x5�5�5�5�5�5�5�5�5�5�5�5666,60646<6T6X6p6�6�6�6�6�6�6�6�6�6�6�6�6�6�67$7(7,70787P7T7l7p7�7�7�7�7�7�7�7�7�7�7�7�7 88888$8<8L8P8`8d8h8l8p8x8�8�8�8�8�8�8�8�8�8�8 999$94989H9L9P9T9\9t9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 ::(:,:<:@:D:H:L:P:X:p:�:�:�:�:�:�:�:�:�:�:�: ;;;;;,;<;@;P;T;\;t;�;�;�;�;�;�;�;�;�;�;�;�;�; << <0<4<D<H<P<h<x<|<�<�<�<�<�<�<�<�<�<�<�<�<===(=,=4=L=\=`=p=t=�=�=�=�=�=�=�=�=�=�=�=>>>>$><>L>P>`>d>h>p>�>�>�>�>�>�>�>�>�>�>�>�> ???$?4?8?H?L?P?X?p?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? � �  0 0$04080@0X0h0l0|0�0�0�0�0�0�0�0�0�0�0�0�01�1�1�1�1�1�1�1�1�1�1�1�1�1�1�122,242H2P2X2`2d2t2�2�2�2�2�2�2 3333(383\3h3p3�3�3�3�3�344 4@4d4p4x4�4�4�4�4�45 5(5H5l5x5�5�5�5�5�5�56(606P6t6�6�6�6�6�6�6 7$70787X7|7�7�7�7�7�7�78,888@8X8d8�8�8�8�8�8�8�8�8�8�8�8999 9$9(909D9`9�9�9�9�9�9:(:H:h:�:�:�:�:�:�: ; ;@;`;�;�;�;�;�;<<0<P<p<�<�<�<�<�<�<�<=,=8=@=p=x=|=�=�=�=�=�=�=�=�=�=�=>>,>0>P>p>�>�>�>�>?,?0?P?p?|?�?�?�?   � $   0040P0l0�0�0�0�01$1`1�1�1�1�182�2�2�283T3�3�3�3�3404L4h4�4�4�4�4�45D5p5�5�5�5�5�5�5�5�5�5�5�6�6�6H9L9P9�=�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   � �   X0h0x0�0�0�0�0�0�0�0�0�0�0`2d2h2l2p2t2x2|2�2�2�384<4@4D4H4L4P4T4X4\4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5l6t6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67777$7,747<7D7L7�7�7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        