MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��u=��n��n��n��n��n���n��n���n �n�;`n��n��n��n���n��n���n��n���n��nRich��n                        PE  L �4LM        � !	  �  �      .     �                         �                              ` R   � <                            ` �8  ��                            �� @            � \                          .text   ݂     �                   `.rdata  �w   �  x   �             @  @.data   L;                       @  �.reloc  �D   `  F                @  B                                                                                                                                                                                                                                                                                                                                                                                        U�존=V��H�Q`V�ҡ�=�U�H�E�IdRj�PV�у���^]� ���������̡�=�P�BlQ��Y�U��j�hpd�    PQV�'3�P�E�d�    ��u��L �N�E�    ���M> �N$�E��q� �ƋM�d�    Y^��]����������������U��j�hApd�    PQV�'3�P�E�d�    ��u����N$�E�   �¯ �N�E� �f> ���E������(L �M�d�    Y^��]���������U���T  �'3ŉE�Wj j�W= ����u_�M�3���� ��]�V������PWǅ����(  �$= ����   ������Qj�= �����   ������RPǅ����$  ��< ���}   ������P������h  Q�� ������h  R�� ���������P�I �@��u�+�$    ��/t��t������H��\uꍴ����V��� h�V�� ����u.������PW�P< ���8���W� �^3�_�M�3���� ��]ËM�^3͸   _�� ��]���������j j j��l �����U��j�h�pd�    P��`SVW�'3�P�E�d�    ��E�P�M�Q3ۋ��E�   �]���T 9]��2  �M��*� ��=�B�P`�M�Q�]��҃��E�Pj�M܍~Q���E��j@ P�M��E��=� �U�R�M��E��=� �M��E�聭 ��=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�]��у�h���M�跬 �U�R�M��E��� �M��]��,� �E�SP�� �����X  ��=�Q�J`�E�P�ы�=�B�PdSj��M�h��Q�ҍE�P�E�� ��=�Q�Jl�E�P�]��у�S���NL ��=�B�P`�M�Q�ҡ�=�H�AdSj��U�hx�R�ЍM�jQ�E��� ��=���B�Pl�M�Q�E�]��҃� S8]���   hh��M������E�P�E��� ��=�Q�Jl�E�P�]������ h�h�   h�=h�   �E��K� ���E��E�;�t	���ƚ  �3��U�WR�Ȉ]���  h�  ���gK �S�E�P���E�   �]��� �M��E�����谫 �M�d�    Y_^[��]� ������������U���SVW��j�~W�E�3�P�E�   �]��:� jW�M�Q���E�   �]��"� jW�U�R���E�   �]��ZT jW�E�P���E�   �]���S jW�M�Q���E�   �]���S jW�U�R���E�   �]��S j
W�E�P���E�
   �]���S j	W�M�Q���E�	   �]��S jW�U�R���E�   �]��jS j�E�   �]�W�E�P���RS jW�M�Q���E�   �]��J� jW�U�R���E�   �]��"S _^[��]������������U��j�h�qd�    P���   SVW�'3�P�E�d�    ���o ����   h���M��y� ��l���3�P�]��� �M�QP�U�R�E��� ���~$P���E��ī �M��E��ȩ ��l����]�躩 �M��E�����諩 �^@�� �E�SW�E�   �� ������  �E�P���L� P�M��E��� Sj�M�Q�M��E��� ���M��E��E��J� ��=�B�Pl�M�Q�E��҃�8]�t'�E�P�E������,� ��3��M�d�    Y_^[��]�Sh���M��7����M�Q�~j���E��c> ��=�B�Pl�M�Q�E��҃�h��M��-� h���l����E��� ��4���j	P�E��� ��l���QP��P���R�E�	蟪 �M�QP�U�R�E�
荪 �� ��P����E��[� ��4����E��L� ��l����E��=� �M��E��1� �E�jP�� ���M���tQ�M��� Pj���E��= �M��OSh���5���P�E�� ��=�H�Al�U�R�E��Ѓ�Sh���M������M�Qj���E��4= �M܋�=�B�PlQ�E��҃�Sj���< jj����; jj����; jj����; Sj
����; jj	���; jj���; Sj���; Sh���M��x����E�Pj���E��< ��=�Q�Jl�E�P�E��у�Sj���T; �M�W�[� �M��c� �M��E��� �U�R�N$諧 P�M��E��n� �M�Sj�E�P�E���� ���M��E��E�試 ��=�Q�Jl�E�P�E��у�8]�t'�U�R�E������� ��3��M�d�    Y_^[��]ËM�j�~W�F� �M��� ��=�E�   �]�H�A`�U�R�Ѓ��M�Qj�U�R���E���8 SSP�E�P���E��J ��=�Q�Jl�E�P�E��ы�=�B�Pl�M�Q�E��ҡ�=�E�   �]�H�A`�U�R�Ѓ��M�Qj�U�R���E��j8 SSP�E�P���E��8J ��=�Q�Jl�E��E�P�ы�=�B�Pl�M�Q�E��҃�h���h  �Sjh���h  �Sj���E�   �]��6 P�E�P���F SSj���E�   �]��]6 P�M�Q���a� SSj���E�   �]��<6 P�U�R���@� SSj���E�   �]��6 P�E�P���� h���h  �Sjh���h  �Sj
���E�
   �]��6 P�M�Q���F �E�	   �]�SSj	����5 P�U�R���Ǎ SSj���E�   �]��5 P�E�P��覍 SSj���E�   �]��5 P�M�Q��腍 ��=�E�   �]�B�P`�M�Q�҃��E�Pj�M�Q���E���6 SSP�U�R���E��H ��=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��у�SS�E�   �]�j����4 P�U�R����� h�  ���$C �E�P�E�����蔽 ���   �M�d�    Y_^[��]�����������U��j�h�qd�    P��0VW�'3�P�E�d�    ���@ ��   �(� �E��E�P�O$�E�    �� P�M��E�襢 j j�M�Q�M��E��1� �Mċ��E��� ��=�B�Pl�M�Q�E� �҃���t���/����M���W�� �M��� �E�P�E�����諼 ���M�d�    Y_^��]��������U��j�hlrd�    P��   SVW�'3�P�E�d�    ��3ۉ]��F@   �����E����   ����   ���  ��=�H�A`�U�R�Ћ�=�Q�JdSj��E�hh�P�эU�R�E�   �� ��=�H�Al�U�R�E��������l� h�h�   h�=h�   ����� ��,�E�E�   ;�t	���i�  �3���VW���E�����貿  �p  �MQ�U�R���E�   �]��tH 9]�N  h�  ����@ �=  ��� h�h�   h�=j$���m� ��;�t�@   ��X�X�X�X�3���VW���E�������F  ��=�H�A`�U�R�Ѓ��M�Qj�Uؿ   R�Ή}��3 ��=�H�Al�U�R�E��Ѓ�Sj����1 ��t7Sh���M��������=�Q�R S�E�P�M�Q�E��}��҃��E��u�]�E��E�   t��=�H�Al�U�R�Ѓ�8]�  ����S����   ��=�Q�JP�E�P�ы�=���B��H  h��h�   V�ы�=S���B�PTV�M�WQ��j<��L���SP��� ��0��L���QǅL���<   ��P�����T���ǅX���4���\�����d���ǅh���   ��l����T���ueSh��M������U�R�E��"� ��=�H�Al�U�R�E����0h��M������M�Q�E���� ��=�B�Pl�M�Q�E��҃���=�H�Al�U�R�E������Ѓ��   �M�d�    Y_^[��]� ����V��V��� ���    ^�������������VW��3�9>t	V� � ���>�~�~�~�~_^�������������U��V�������Et	V�	� ����^]� �������������������������������U�존=�UV��H�ApVR�Ѓ���^]� ��������������U�존=V��H�Q`V�ҡ�=�H�U�ApVR�Ѓ���^]� ��=���   �Q��Y���������������U������P�M�P��P�P�P�P �P�P�P,�P(�X$���Q�P�I�H�M��P�Q�P�I�H�M��P�Q�P�I�H �M��P$�Q�P(�I�H,]� ���U��M�U�A�
�E��A�J���A$�J����A�
�A�A�J���A(�J���X�A�
�A�A �J���A,�J���X�A�J�A�J���B�I$���X�A�J�A�J���B�I(���X�A �J�A�J���A,�J���X�A�J�A�J���B �I$���X�A�J�A�J���B �I(���X�A �J�A�J���A,�J ���X �B$�I�A�J(���B,�I$���X$�A�J(�A�J$���B,�I(���X(�A �J(�A�J$���A,�J,���X,]���U��j�h�rd�    P��SVW�'3�P�E�d�    3ۉ]�]��E�M�Q�M�]��E؉]܉]��� �}S�U�R�E�P���E��! �M���]��a ;�t}��=���   �JX�E�P�ы���;�t_��=���   �PT���ҋ�=���   �M�RQPV�ҋ�=���   ��U�R�E������Ѓ��ƋM�d�    Y_^[��]� ��=���   �
�E�P�E������у�3��M�d�    Y_^[��]� ������������U��j�h�rd�    P�� SVW�'3�P�E�d�    3ۉ]��]�]�E�M�Q�   �M��}��Eԉ]؉]�� �MS�U�R�E�P�E��  �M����E��* ;�t\��=���   �JH�E�P�ы�=�u���B�H`V�ы�=�B�HpVW�ы�=���   ��M�Q�E�   �]��҃��C��=�H�u�Q`V�ҡ�=�H�QdSj�h��V�ҡ�=���   ��U�R�}��]��Ѓ��ƋM�d�    Y_^[��]� �U��j�hsd�    P��SV�'3�P�E�d�    3ۉ]�]��E�M�Q�M�]��E؉]܉]�� �MS�U�R�E�P�E��a �M���]�� ;�tJ��=���   �J8�E�P�ы�=�����   ��M�Q�E������҃��ƋM�d�    Y^[��]� ��=���   ��U�R�E������Ѓ�3��M�d�    Y^[��]� ����U��j�hKsd�    P�� SV�'3�P�E�d�    3��u��u�u�E�M�Q�M��u��Eԉu؉u�� �MV�U�R�E�   P�]��]��g ��t��=���   �J�E�P�у���u2ۍM��u���	 ��tK��=���   �P<�M�Q���]��=���   ��U�R�E��������E���M�d�    Y^[��]� ��=���   �
�E�P�E��������E���M�d�    Y^[��]� �������U��j�hvsd�    P��SV�'3�P�E�d�    3ۉ]�]��E�M�Q�M�]��E؉]܉]�� �MS�U�R�E�P�E��Q �M���]��� ��=���   �E�P;�t7�J@�ы�u�H��P��=�N���   ��V�U�R�E������Ѓ����u�
�V�V�E�������у��ƋM�d�    Y^[��]� ���������U��j�h�sd�    P�� SV�'3�P�E�d�    3ۉ]��]�]�E�M�Q�M��E�   �Eԉ]؉]�� �MS�U�R�E�P�E��Z �M����E��� ;�tC��=���   �JL�E�P�ыu��P����� ��=���   ��M�Q�E�   �]����(�uS���j� ��=���   ��U�R�E�   �]��Ћƃ��M�d�    Y^[��]� �����U��j�h�sd�    PQSVW�'3�P�E�d�    ��=�H�AP�Uj3�R�}��Ћ�=�Q����H  h@�Fh�  V�Ћ�=j�E��Q�JTVP�EP��N��$;�~�]�U��P����� G;�|�M�Q�� ��=�B�Pl�MQ�E������҃��M�d�    Y_^[��]� ��U��j�h td�    P��SVW�'3�P�E�d�    ��=�H�A`�U�R�Ћ�=�Q�Jd3�Wj��E�h��P�ы�=�B�PP�M�jQ�}��ҋ�=�H��H  h@�Fh�  V�ҋ�=j�E��Q�JTVP�E�P��N��8;�~�]���U��P����� G;�|�M�Q�� ��=�B�Pl�M�Q�E������҃��M�d�    Y_^[��]� ���U��Q�ESVW���   3�3�3�3ۃ��M�|#�@|�O���A�	�d$ p����u�E�M�;�}�@|��_�^�[��]� �����U��j�h�td�    P��   SV�'3�P�E�d�    3ۉ]�=�H�u�Q`V�]��ҡ�=�H�QdSj�h0�V�҃��E�]��E�   ��
�j  �$��0 Sh,��M��I����E�P���E�   �W_  ��=�Q�Jl�E�P�]����&  Sh(��M������U�R���E�   �_  �U���  Sh ��M�������M�Q���E�   ��^  ��=�B�Pl�M�Q�]�����  Sh���p���������p���P���E�   �^  ��=�Q�Jl��p���P�]����  Sh��M��j����U�R���E�   �x^  �U��H  Sh���P����?�����P���Q���E�   �J^  ��=�B�Pl��P���Q�]����  Sh��M�������E�P���E�   �^  ��=�Q�Jl�E�P�]�����   Sh��M�������U�R���E�   ��]  �U��   Sh���M������M�Q���E�	   �]  ��=�B�Pl�M�Q�]����}Sh����`����c�����`���P���E�
   �n]  ��=�Q�Jl��`���P�]����=Sh���@����#�����@���R���E�   �.]  ��@�����=�H�AlR�]��Ѓ���=�Q�J`�E�P�ы�=�B�PdSj��M�h�Q�ҡ�=�H�QV�E�   �ҋ�=�Q�R0�M�QPV�ҡ�=�H�Al�U�R�]��Ѓ�(�ƋM�d�    Y^[��]� �I �- �- . E. �. �. �. -/ U/ �/ �/ ����U��j�hud�    PQSVW�'3�P�E�d�    ���}�3��   �G�7�w�w�w�w�_�u��C�3�s�s�s�s�G@�w0�w4�wD�w<�w8�GX�wH�wL�w\�wT�wP�Gp�w`�wd�wt�wl�wh���   �wx�w|���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   ���   �E�97t	W�\� ���7�w�w�w�w93t	S�A� ���G0�3�s�s�s�s90t	P�#� ���GH�w0�w4�wD�w<�w890t	P�� ���G`�wH�wL�w\�wT�wP90t	P�� ���Gx�w`�wd�wt�wl�wh90t	P�ƺ �����   �wx�w|���   ���   ���   90t	P蛺 �����   ���   ���   ���   ���   ���   90t	P�j� �����   ���   ���   ���   ���   ���   �ǋM�d�    Y_^[��]����������������U��j�h�ud�    PQSVW�'3�P�E�d�    ��u��E�   ��� ���   3��E�9t	W�ӹ ����_�_�_�_���   �E�9t	W讹 ����_�_�_�_�~x�E�9t	W茹 ����_�_�_�_�~`�E�9t	W�j� ����_�_�_�_�~H�E�9t	W�H� ����_�_�_�_�~0�E�9t	W�&� ����_�_�_�_�~�]�9t	W�� ����_�_�_�_�E�����9t	V�� ����^�^�^�^�M�d�    Y_^[��]�U��j�h�vd�    P��(  SVW�'3�P�E�d�    ���}존=�H�A`�U�R�Ћ�=�Q�Jdj j��E�hP�P�ы�=�B�P`��|���Q�E�    �ҡ�=�H�Adj j���|���hD�R�ЋMQ�����R�E�� P��|���P��<���Q�E��X  �U�RP�E�P�E��X  ��H��=�Q�Jl��<���P�E��ы�=�B�Pl�����Q�E��ҡ�=�H�Al��|���R�E��Ћ�=�Q�Jl�E�P�E��ы]��=�B�H`��S����e�V�ы�=�B�Pp�M�VQ�҃����/����u�~ �E�    �e  3���=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�ы�=�B�P`�M�Q�E�	�ҡ�=�H�Adj j��U�h@�R�Ћ�=�Q�J`��\���P�E�
�ы�=�B�Pdj j���\���h@�Q�ҡ�=�H�A`�U�R�E��Ћ�=�Q�Jd��@j j��E�h<�P�у��F�D8j0j jj �Q�U��$�E�R�~ ���؋F�D8j0j j�j Q��L����$P�E��T ���E�F�8j0j j�j Q��l����$Q�E��* P�U�R��,���P�E��V  ��\���QP������R�E��}V  �MQP������R�E��hV  �M�QP�����R�E��SV  ��HSP������P�E��>V  �M�QP������R�E��)V  ��=�Q�Rp�M�QP�E��ҡ�=�H�Al������R�E��Ћ�=�Q�Jl������P�E��ы�=�B�Pl�����Q�E��ҡ�=�H�Al������R�E��Ћ�=�Q�Jl������P�E��ы�=�B�Pl��,���Q�E��ҡ�=�H�Al��l���R�E��Ћ�=�Q�Jl��L���P�E��ы�=�B�Pl�M���@Q�E��ҡ�=�H�Al�U�R�E����E�
��=�Q�Jl��\���P�ы�=�B�Pl�M�Q�E�	�ҡ�=�H�Al�U�R�E��ЋM��=�B��Q�H`���܉eS�ы�=�B�Pp�M�SQ�ҋM��������E�@��;F�E�������}�]��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�hP�P�ы�=�B�P`�M�Q�E��ҡ�=�H�Adj j��U�h4�R�ЋMQ��l���R�E��� P�E�P��L���Q�E��T  �U�RP�E�P�E���S  ��H��=�Q�Rp�M�QP�E��ҡ�=�H�Al�U�R�E��Ћ�=�Q�Jl��L���P�E��ы�=�E��B�Pl��l���Q�ҡ�=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��ы�=�B�H`��S����eV�ы�=�B�Pp�M�VQ�҃����[���S���#�����=�H�Al�U�R�E������Ѓ��M�d�    Y_^[��]� ����U��j�h<yd�    P��  SVW�'3�P�E�d�    ���}衴=�H�A`������R�Ћ�=�Q�Jdj j�������hl�P�ы�=�B�P`�����Q�E�    �ҡ�=�H�Adj j������hD�R�Ћu�F,P������Q�E�� P�����R��(���P�E��&R  ������QP�U�R�E��R  ��H��=�H�Al��(���R�E��Ћ�=�Q�Jl������P�E��ы�=�B�Pl������E�Q�ҡ�=�H�Al������R�E��ЋM��=�B��Q�H`���܉eS�ы�=�B�Pp�M�SQ�҃�������3�9]�]�  ��=�H�A`������R�Ћ�=�Q�Jdj j�������h��P�ы�=�B�P`��x���Q�E�	�ҡ�=�H�Adj j���x���h@�R�Ћ�=�Q�J`������P�E�
�ы�=�B�Pdj j�������h@�Q�ҡ�=�H�A`������R�E��Ћ�=�Q�Jd��@j j�������hh�P�у��Fj0�<[j �j��D8�j �E�Q��(����$R�� ���E��F�D8���j0j ��jj Q�]썅����E��E��$P� ���E�F�8j0j j�j Q�������$Q�E��} P������R��x���P�E���O  ������QP��H���R�E���O  �M�QP��H���R�E��O  ��x���QP��h���R�E��O  ��H�M�QP��X���R�E��O  ������QP��x���R�E��pO  ��=�Q�Rp�M�QP�E��ҡ�=�H�Al��x���R�E��Ћ�=�Q�Jl��X���P�E��ы�=�B�Pl��h���Q�E��ҡ�=�H�Al��H���R�E��Ћ�=�Q�Jl��H���P�E��ы�=�B�Pl��x���Q�E��ҡ�=�H�Al������R�E��Ћ�=�Q�Jl�����P�E��ы�=�B�Pl��@��(���Q�E��ҡ�=�H�Al������R�E��Ћ�=�Q�Jl������P�E�
�ы�=�B�Pl��x���Q�E�	�ҡ�=�H�Al������R�E��ЋM��=��Q�J�Q`���ĉe�P�E��ҡ�=�H�U��IpR�E�P�ыM��������=�B�P`������Q�ҡ�=�H�Adj j�������h��R�Ћ�=�Q�J`�E�P�E��ы�=�Bj j�h@��M�Q�Pd�ҡ�=�H�A`������R�E��Ћ�=�Q�Jdj j�������h@�P�ы�=�B�P`��X���Q�E��ҡ�=�H�Ad��@j j���X���hh�R�Ѓ��N�Dj0j j�Dj Q��h����$R�E��Y
 ���E�F�D�D��j0j ��jj Q�]��������E��E��$Q�"
 ���E��Vj0j �E��|j�j Q�������$P��	 P��X���Q������R�E��_L  ������QP������R�E��GL  �M�QP�����R�E��2L  �M�QP������R�E��L  ��H�M�QP������R�E� �L  ������QP������R�E�!��K  ��=�Q�Rp�M�QP�E�"�ҡ�=�H�Al������R�E�!�Ћ�=�Q�Jl������P�E� �ы�=�E��B�Pl������Q�ҡ�=�H�Al�����R�E��Ћ�=�Q�Jl������P�E��ы�=�B�Pl������Q�E��ҡ�=�H�Al������R�E��Ћ�=�Q�Jl������P�E��ы�=�B�Pl��h�����@Q�E��ҡ�=�H�Al��X���R�E��Ћ�=�Q�Jl������P�E��ы�=�B�Pl�M�Q�E��ҡ�=�H�Al������R�E��ЋM��Q���e���=�B�H`��W�ы�=�B�Pp�M�WQ�ҋM��������=�H�A`��h���R�Ћ�=�Q�Jdj j���h���h��P�ы�=�B�P`�M�Q�E�#�ҡ�=�H�Adj j��U�h@�R�Ћ�=�Q�J`�E�P�E�$�ы�=�B�Pdj j��M�h@�Q�ҡ�=�H�A`�����R�E�%�Ћ�=�Q��@j j�hh������P�Jd�у��Fj0j �|[�j��D8�j Q��x����$R�E�&�� ���E�F�D8���j0j ��jj Q�]��������E��E�'�$P� ���E��F�8j0j j�j Q�������$Q�E�(� P�����R������P�E�)��H  �M�QP������R�E�*��H  �M�QP�����R�E�+�H  �M�QP��8���R�E�,�H  ��H�M�QP��X���R�E�-�H  ��h���QP��h���R�E�.�xH  ��=�Q�Rp�M�QP�E�/�ҡ�=�H�Al��h���R�E�.�Ћ�=�Q�Jl��X���P�E�-�ы�=�B�Pl��8���Q�E�,�ҡ�=�H�Al�����R�E�+�Ћ�=�Q�Jl������P�E�*�ы�=�B�Pl������Q�E�)�ҡ�=�H�Al�������E�(R�Ћ�=�Q�Jl������P�E�'�ы�=�B�Pl��x�����@Q�E�&�ҡ�=�H�Al�����R�E�%�Ћ�=�Q�Jl�E�P�E�$�ы�=�B�Pl�M�Q�E�#�ҡ�=�H�Al��h���R�E��ЋM��=�B��Q�H`�����e�W�ы�=�B�Pp�M�WQ�ҋM�������N|�E�<��u  ��=�B�P`�M�Q�ҡ�=�H�Adj j��U�h��R�Ћ�=�Q�J`�E�P�E�0�ы�=�B�Pdj j��M�h@�Q�ҡ�=�H�A`��(���R�E�1�Ћ�=�Q�Jdj j���(���h@�P�ы�=�B�P`��H���Q�E�2�ҡ�=�H�Ad��@j j���H���hh�R�Ѓ��Fj0�|[	j �j��D8�j �E�3Q��8����$Q�\ ���E�F�D8���j0j ��jj Q�]��������E��E�4�$R�' ���E��F�8j0j j�j Q�������$P�E�5�� P��H���Q������R�E�6�eE  ��(���QP������R�E�7�ME  �M�QP������R�E�8�8E  �M�QP�����R�E�9�#E  ��H�M�QP��8���R�E�:�E  �M�QP��X���R�E�;��D  ��=�Q�Rp�M�QP�E�<�ҡ�=�H�Al��X���R�E�;�Ћ�=�Q�Jl��8���P�E�:�ы�=�B�Pl�����Q�E�9�ҡ�=�H�Al������R�E�8�Ћ�=�Q�Jl������P�E�7�ы�=�B�Pl������Q�E�6�ҡ�=�H�Al������R�E�5�Ћ�=�Q�Jl������P�E�4�ы�=�B�Pl��@��8���Q�E�3�ҡ�=�H�Al��H���R�E�2�Ћ�=�Q�Jl��(���P�E�1�ы�=�B�Pl�M�Q�E�0�ҡ�=�H�Al�U�R�E��ЋM��=�B��Q�H`�����e�W�ы�=�B�Pp�M�WQ�ҋM�������E�N|�@;E�E������}��=�B�P`�M�Q�ҡ�=�H�Adj j��U�hl�R�Ћ�=�Q�J`�E�P�E�=�ы�=�B�Pdj j��M�h4�Q�ҋv,������VP�E�>�� P�M�Q������R�E�?��B  �M�QP��8����@R�]��B  ��H��=�Q�Rp�M�QP�E�A�ҡ�=�H�Al��8���R�]��Ћ�=�Q�Jl������P�E�?���E�>��=�B�Pl������Q�ҡ�=�H�Al�U�R�E�=�Ћ�=�Q�Jl�E�P�E��ы]��=�B�H`��S����eV�ы�=�B�Pp�M�VQ�҃�������S���������=�H�Al�U�R�E������Ѓ��M�d�    Y_^[��]� �U��j�h�zd�    P���   SVW�'3�P�E�d�    ��=�HH�U���  j h�  R�Ћ}��j j�ωE�� j j�ωE��v ��=�Q�J`���E�P�}��у��E�    ���4  �~ �*  ��\����Hs ��0���R�E�舾 ���!� P��\����E��u ��0����E���s ��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�у��U�R��\����E���t ��=�H�Al�U�R�E��Ћ�=�Q�J`�E�P�ы�=�B�Pdj j��M�h��Q�ҡ�=�H�A`�U�R�E��Ћ�=�Q�Jdj j��E�h��P�у�,�E���0���R��\����E� �M�Q���E��s P�U�R�E�P�E���?  �M�QP�U��R�]���?  ��=�Q�Rp�M�QP�E�	�ҡ�=�H�Al�U�R�]��Ћ�=�Q�Jl�E�P�E��ы�=�B�Pl�M�Q�E��҃�,��0����E��Xr ��=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��ы]��S���e����=�B�H`W�ы�=�B�Pp�M�WQ�҃����2���S���������\����E� ��q ��]��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�ы�=�B�P`�M�Q�E�
�ҡ�=�H�Adj j��U�h��R�Ѓ�(��=���   �M�Bx�E���P�M�Q�U�R�a>  �M�QP�U�R�E��O>  ��=�Q�Rp�M�QP�E��ҡ�=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��ы�=�B�E�
�MċPlQ�ҡ�=�H�Al�U�R�E� �Ћ�=�Q�B`��0S�����eW�Ћ�=�Q�Jp�E�WP�у��������S�������U�}RWS���"����}� t�E��MPQWS��������=�B�P`�M�Q�ҡ�=�H�Adj j��U�h��R�Ћ�=�Q�J`�E�P�E��ы�=�B�Pdj j��M�hD�Q�ҋEP�M�Q�E���� P�U�R�E�P�E���<  �M�QP�U�R�E���<  ��H��=�Q�Rp�M�QP�E��ҡ�=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��ы�=�E��B�Pl�M�Q�ҡ�=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E� �ы�=�J�Q`��S���ĉeP�E�ҡ�=�H�U�IpR�E�P�у����V�����=�B�P`��L���Q�E    �ҡ�=�H�Adj j���L���h��R�Ћ�=�Q�J`��x���P�E��ы�=�B�Pdj j���x���h��Q�҃�(�} �E��E    �  �}� ��  �~ ��  ���   �M�������   ��=��� ���   �ȋBx�Ћ�=�Q�Rp��x���QP�ҡ�=�H�I j ��L���R��x���P�у����_  ��=�B�P`�M�Q�ҡ�=�H�Adj j��U�h��R�Ћ�=�Q�J`�E�P�E��ы�=�B�Pdj j��M�h��Q�ҍ�x���P�M�Q�� ���R�E��:  �M�QP�� ���R�E��:  ��@��=�Q�Rp�M�QP�E��ҡ�=�H�Al�� ���R�E��Ћ�=�Q�Jl�� ���P�E��ы�=�B�Pl�M�Q�E����E���=�H�Al�U�R�Ћ�=�Q��S���ĉe�EP�B`�Ћ�=�Q�E�RpP�M�Q�҃���������=�H�Ip��L���R��x���P�у���=�B�P`�����Q�ҡ�=�H�Adj j������h��R�Ћ�=�Q�Rp�E�P�����Q�E��ҡ�=�H�Al�����R�E��ЋO|�U�� �<� �E    ��  �]�����    ��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h@�P�ы�=�B�P�M�Q�E��ҋ�=�Q�M�Q�J0P�E�P�ы�=�B�Pl�M�Q�E��ҋG4�N�ÍDP��<���Q�� �E��=�B�P�M�Q�E��ҋ�=�Q�MQ�J0P�E�P�ы�=�B�Pl��<�����@Q�E��҃��}� ��   �\ ��   ��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�ы�=�B�P�M�Q�E��ҋ�=�Q�M�Q�J0P�E�P�ы�=�B�Pl�M�Q�E��ҋGL�N�ÍDP��h���Q�� �E��=�B�P�M�Q�E��ҋ�=�Q�MQ�J0P�E�P�ы�=�B�Pl��h�����@Q�E��҃��E�O|�U@��;��E�����]��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�ы�=�B�P�M�Q�E��ҋ�=�Q�M�Q�J0P�E�P�ы�=�B�Pl�M�Q�E��ҋ�=�Q��(S���ĉe�EP�B`�Ћ�=�Q�E�RpP�M�Q�҃���������E�O|��U@;E�E�������=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�ы�=�B�P`�M�Q�E��ҡ�=�H�Adj j��U�h4�R�ЋMQ�� ���R�E� ��� P�E�P��<���Q�E�!�6  �U�RP��h���P�E�"��5  ��H��=�Q�Rp�M�QP�E�#�ҡ�=�H�Al��h���R�E�"�Ћ�=�Q�Jl��<���P�E�!�ы�=�E� �B�Pl�� ���Q�ҡ�=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��ы�=�B�H`��S�����eW�ы�=�B�Pp�M�WQ�҃����U���S��������=�H�Al��x���R�E��Ћ�=�Q�Jl��L���P�E� �ы�=�B�Pl�M�Q�E������҃��M�d�    Y_^[��]� ������������U��j�h�{d�    P��  SVW�'3�P�E�d�    ��=�H�A`��`���R�E�    �Ћ�=�Q�Jdj j���`���h@�P�э�`���R�EP�M�Q�E��24  ��=�B�Pl��`���Q�E��ҋE�]��$PS�M�Q���C�����=�B�P`�M�Q�ҡ�=�H�Adj j��U�h��R�Ћ�=�Q�J`�E�P�E��ы�=�B�Pdj j��M�h@�Q�ҡ�=�H�E���p����A`R�Ћ�=�Q�Jdj j���p���h@�P�у�<�E�j0j jj Q�U��$R�E���� �����E�j0j jj Q�E��$P�E��� ���E�E�j0j jj Q��P����$Q�E��� ��p���RP��4���P�E�	��2  �MQP�����R�E�
��2  �M�QP������R�E���2  W�E�P������P�2  ��H�M�QP�����R�E��2  ����=�H�A�U�R�E��Ћ�=�Q�J0WP�E�P�ы�=�B�Pl�����Q�E��ҡ�=�H�Al������R�E��Ћ�=�Q�Jl������P�E��ы�=�B�Pl�����Q�E�
�ҡ�=�H�Al��4���R�E�	�Ћ�=�Q�Jl��P���P�E��ы�=�B�Pl�M�Q�E��ҡ�=�H�E��Al�U�R�Ћ�=�Q�Jl��p���P�E��ы�=�B�Pl�Mă�@Q�E��ҡ�=�H�Al�U�R�E��ЋM��=�B��Q�H`�����eW�ы�=�B�Pp�M�WQ�҃����c����Eh�  PS����������~  h�  P��(���Q���6�����D����E��7c ��M��]��*c ���M�U�R�E��Ƞ ��D���QW��(���RP�E��_� ���M��E��c �M��]��c ��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h@�P�ы�=�B�P`�M�Q�E��ҡ�=�H�Adj j��U�h��R�ЍMQ�U�R�E�P�E��40  �E��M�QP�U�R�"0  ��@��=�Q�Rp�M�QP�E��ҡ�=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��ы�=�B�Pl�M�Q�E��ҡ�=�H�Al�U�R�]��Ћ�=�Q�J`�E�P�ы�=�B�Pdj j��M�h��Q�҃�,�E�P��D����E��0c �M�QP�U�R�E��^/  ����=�H�U��E�R�A�Ћ�=�Q�J0WP�E�P�ы�=�B�Pl�M�Q�E��ҡ�=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�]��ыU��=�H��(R�Q`�����eW�ҡ�=�H�Ap�U�WR�Ѓ����������D����E��a ��(����E��a ��=�Q�Jl�E�P�E� �ы�=�B�Pl�MQ�E������҃��M�d�    Y_^[��]�$ ������U��j�h]|d�    P���   SVW�'3�P�E�d�    ��M��[` ��=�H�A`�U�R�E�    �Ѓ��M�Q�M�   S�U�R�E���  P��D����]��g` ��D���P�M��E��db ��D����]��` ��=�Q�Jl�E�P�E��ы�=�B�Pl�M�Q�E� �ҋM����D���P訜 P�M��E��+b ��D����E� �L` ��=�Q�J`�E�P�ы�=�B�Pdj j��M�h��Q�҃��E��E�P�M��|a ��=�Q�Jl�E�P�E� �у��U�R�M��` P�E�荹 ��=�H�Al�U�R�E� �Ѓ��c �E�h1D4ChCD4C�E����(� Pj S�M�Q���c ��u;�U�R�E��Yc ���M��E�    �E������p_ 3��M�d�    Y_^[��]� �~ �E    ��  �F�M��=�<��B�P`�M�Q�ҡ�=�H�A`��p���R�E��Ћ�=�Q�Jdj j���p���h��P�ы�=�B�P`�M�Q�E�	�ҡ�=�H�Adj j��U�h�R�Ѓ�,��=���   �Bx���E�
��P�M�Q��P���R�+  ��p���QP��4���R�E��+  ��=�Q�Rp�M�QP�E��ҡ�=�H�Al��4���R�E��Ћ�=�Q�Jl��P���P�E�
�ы�=�B�Pl�M�Q�E�	�ҡ�=�H�Al��p���R�E��ЋM���=�B��0Q�H`���܉e�S�ы�=�B�Pp�M�SQ�҃���������=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h�P�ы�=�B�@p�M�Q�U�R�E��Ћ�=�Q�Jl�E�P�E��ыU�=�� R���e�܋H�Q`S�ҡ�=�H�Ap�U�SR�Ѓ�������h�  W���r�����tL��=�Q�B`���܉e�S�Ћ�=�Q�Bdj j�h�S�ЋM��U��h4  h@  WQR���B���h�  W��������tJ��=�H�Q`���܉e�S�ҡ�=�H�Qdj j�hܤS�ҋE��M��h�	  hD  WPQ���������=�B�P`��`���Q�ҡ�=�H�Adj j���`���h̤R�Ћ�=�Q�Rp�E�P��`���Q�E��ҡ�=�H�Al��`���R�E��ЋM���=�B�� Q�H`�����e�W�ы�=�B�Pp�M�WQ�҃����%�����=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�ы�=�B�@p�M�Q�U�R�E��Ћ�=�Q�E��Jl�E�P�ыU�=�H�� R�Q`�����e�W�ҡ�=�H�Ap�U�WR�Ѓ���������=�Q�J`�E�P�ы�=�B�Pdj j��M�h��Q�ҡ�=�H�Ip�U�R�E�P�E��ы�=�B�Pl�M�Q�E��ҋE���=�Q�� P�B`�����e�W�Ћ�=�Q�Jp�E�WP�у���������U�R��������=�H�Al�U�R�E��ЋE@��;F�E�=����M��^ �M�Q�E� �A^ ���M��E�    �E������XZ �   �M�d�    Y_^[��]� ���������������U��j�h�~d�    P��  SVW�'3�P�E�d�    �ى�����hG  ��� �K ���� ��������  �������"Y ��=�H�A`�U�R�E�    �Ѓ��u�M�Qj�U�R���E��_�  P��(����E��/Y ��(���P�������E��)[ ��(����E��jY ��=�Q�Jl�E�P�E��ы�=�B�Pl�M�Q�E� �ҋ}����(���P���j� P�������E���Z ��(����E� �Y ��=�Q�J`��`���P�ы�=�B�Pdj j���`���h4�Q�҃��E���`���P�������/Z ��=�Q�Jl��`���P�E� �у���������W ��=�B�P`�M�Q�E��҃��E�Pj�M�Q���E��*�  P��(����E���W ��(���R�������E�	��Y ��(����E��5X ��=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��у�h(���(����gW ��(���R�������E�
�Y ��(����E���W �������W ��=�H�U��E�R�A`�Ѓ��M�Qj�U�R���E��Z�  P��(����E��*W ��(���P�������E��$Y ��(����E��eW ��=�Q�Jl�E�P�E��ы�=�B�Pl�M�Q�E��҃�h���(����V ��(���P�������E���X ��(����E��W �M�Q��������W P�E�蘰 ��=�B�Pl�M�Q�E��҃��E�P�������W P�E��f� ��=�Q�E��E؋JlP�у��U�R�������^W P�E��4� ��=�H�Al�U�R�E������Ũ��UЍM���Q�]ԍ����R��H���ٕ���P�荍d���ٕ ���QٝH�����x���ٕ$���ٕL���ٕP���ٕd���ٕh���ٝl���������=���   ���   �щE�j P���E�芎 ��=���   �M苐�   �҅���  �vY �E�h1D4ChCD4C�E����� Pj j������P���Y ��uz�M�Q�E��JY ��=3��u싂�   ���   �M�Q�E��҃��u荍�����E��DU �������E� �5U �������E������#U 3��M�d�    Y_^[��]� j h���M��>����E�P�M�Q�������E��U ���ԉečM�QPR�E���!  ����������=�B�Pl�M�Q�E��ҡ�=�H�Al�U�R�E��Ѓ�j h���M��ɣ���M�Q�U�R�������E��BU ���̉ečU�RPQ�E��k!  ����葾����=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��у�j h���M��T����U�Rj j���E��q�  P�E�P���e������̉ečU�RPQ�E���   ����������=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��у�j j����  P�U�R�������P�E��5� ��=�H�Al�U�R�E��ЋM���W j h��M�薢��j h ��M��E�胢��������E�Q��������S P�U�R��`���P�E��(   �M�QP�����R�E��   P�E� 詬 ��=�H�Al�����R�E��Ћ�=�Q�Jl��`���P�E��ы�=�B�Pl�����Q�E��ҡ�=�H�Al�U�R�E��Ћ�=�Q�Jl�E�P�E��у�0�<V �E�h1D4ChCD4C�E�!���� Pj j������R���QV ��u6�E�P�E��V �M�3�Q�u��E���U ���M�u��E���  �������=�B�P`��D���Q�҃�3�Whܥ�M��E�"�+�����=�H�Ip��D���R�E�P�E�#�ы�=�B�Pl�M�Q�E�"�ҋE���P����D����̉e�R�n������׻���   ��4�����0�����,���Pǅ,����  ��@�����<�����8����n ��Wh���M�荠��Wh̥�M��E�$�{�����,���Q�����h��R�E�%�O P�E�P��`���Q�E�&�  �E�'�U�RP�����P�  ��$P��D����E�(育����=�Q�Jl�����P�E�'�ы�=�B�Pl��`���Q�E�&�ҡ�=�H�Al�����R�E�%�Ћ�=�Q�Jl�E�P�E�$�ы�=�B�Pl�M�Q�E�"�ҋE���P����D����̉e�R�!�����芺��Wh���M��|���Wh���M��E�)�j�����=� P�����Q�E�*�� P�U��E�+R��`���P�  �M�QP�����R�E�,��  �� P��D����E�-�u�����=�H�Al�����R�E�,�Ћ�=�Q�Jl��`���P�E�+�ы�=�B�Pl�����Q�E�*�ҡ�=�H�Al�U�R�E�)�Ћ�=�Q�Jl�E�P�E�"�ыU���R����D����̉e�P�������~����M�Q���C���Wj���i�  �M�{�{��=���������   ���   ��\����҅��z  �C� ��=���   ��\����M苒�   P�ҋ���=���   �B�ω}���=�  �  ��=�Q�J`�����P�ы�=�B�Pdj j������h��Q�҃���=���   �Bx���E�.��P�����Q������R�d  P�E�/�ʨ ��=�H�Al������R�E�.�Ћ�=�Q�Jl�����P�E�"�у�������������=�B�P`�����Q�E�0�ҡ�=�H�Adj j������h��R�Ѓ���=���   �Bx���E�1��P�����Q������R�  P�E�2�M� ��=�H�Al������R�E�1�Ћ�=�Q�Jl�����P�E�0�у������� ��  ��=�BH���   h�  ��V�у�P��p����  j��������  j ��p����J  ���E�    ��� ���u�����  ��=���   �P����=�  ��  hF  h�  V��诰�����{  j ���E�   ��� ������  h�  V�E�P��謱����=�Q�J�E�P�E�7�у�����   W�������_  �M��7� ������   ���$    �d$ ��=���   �P����=)  ��   ��=���   �Bx���ЍM�Q���  ��tu���J� ��X���R������Q3�V�ȉE��/ ��tO�	��$    ��������F;�X������������t���J��@;�X���~�M���X���R������PV�� ��u���=���   �B(���Ћ����/�����������9j ��p����  ��=�B�Pl�M�Q�E�0�ҋu�����=���   �B(���Ћ��E����.����������9 ��   ��=�B�P`�M�Q�ҡ�=�H�Adj j��U�h��R�Ѓ���=���   �� �����@|�U�R�E�8�Ћ�=�Q�Jl�E�P�E�0�ы�=��JT�Q,j P�҃�����
  ������Q���l �荕d���ٕd���Rٕh���h�  ٝl����������E�9��  ���������������E�0���  �}� ��   ������ �E�    ��   ��    3�9{~a���$    �S��=��� ���   �ȋBx�Ћ������Uȋ���=���   �Bx�Ћ�=�Qj VP�B �Ѓ���t1G;{|��s�������Uȋ<���|jjjV����  ��t�C�<��E�@;������E��Z�����=�QH�u����  j h�  V�Ћ�=�QHj ��������  h�  V�Ћ�=�QH�E����   h�  V�Ћ�=�QH�E����   h�  V�Ћ���h�����(�}�;�t(}+�PW��T����  �jj��+�QP��T����  3���~-�u�����I �3�;V��X�����@����;ǉL��|�u��}�������P��蝴����l���������;�t(}+�PW�������  �jj��+�QP�������  ��H���R����� P��x���P��p���Q�Ӫ���E��E����E�3Ƀ��E��E��)  �u����������G����F��    �U�م|����������H�T8��؅p����E��H������H����]̋]��E��H�؅t������H������H����]��E��H�؅x������H������H��]ЉY���]ԋ]�م|����Y�H��������L؅p����E��H���������]̋U��E��H�؅t������H���������]��E��H�؅x������H��������UЉQ���]ԋU�م|����Q�H؅p����E��H������ȍW������H���]̋U��E��H؅t������H�����H���]��E��H؅x������H�����H��UЉQ���]ԋU�م|����Q�H�������W�؅p�����E��H�����H��ٝT����E��H؅t������H�����H���]��E��H؅x������H�����H���]�مT����]̋U��E���]ЋU��E��Q�]ԋUԃ�0���Q������Mċ�����;M���   ������I������D�+�U�+�م|����������H��ȃ���؅p����E��H������H���ٝT����E��H�؅t������H������H����]��E��H�؅x������H������H����]�مT����]̋}��E��9�]Ћ}��E��y�]ԋ}ԉy�f�����l����܋� �����������;�t&}+�QP������  �jj+�PQ������!  3�3�9M�~w�U���X������<������u.�r�4��2������t��r�������t��r�������t���2�4��r�������t��r�������t���X����A��;M�|��Mj j��  ���_  ��=�BH�u��Hxj h'  V�ы�������  ��l��������;�t,}+�QP�������f
  �jj+�PQ�������a  ��l�����8���;�t&}+�QP��$����  �jj+�PQ��$�����  ����� ��ٕx���3�ٕt���3�9u�ٕp����U��E��U��}�ٕ|����U��U��U��U��U��]���  ��=�BD�Uċ@T��p���QWR�Ћ�X����v�����<���   ��������U���U��Q�U��Q�������U��T�D�M��H�U��P�������F�@����|�����U��Q�U��Q�������N�I����p����:��t����z��x����z��(����4���(����V�T���(����}�����(������   �������U���U��T�U��T��|���ȋ������T�D�M��H�U��P�������F�@����p������t����Q��x����Q��(����4���(����V�T���(�������X���4�G;}ȉ}������MȋU��uQ�M�R�U�������PQRV���<���������Cj j����  ��t	�����K�������E�"������=��\������   �M苐�   G��\�����;������3��M��E 9�����t9{~�UVR��������=�H�Al��D���R�E�!�ЍM�Q�E��E �U�R�}��E���D ���|  j h|���`����N���3�Vhd��M��E�3�:�����=���   �M��Bx�E�4��P�M�Q������R��  ��`���QP�������5R�]���  P�E�6�_� ��=�H�Al������R�]��Ћ�=�Q�Jl������P�E�4�ы�=�B�Pl�M�Q�E�3�ҡ�=�H�Al��`���R�E�0�Ѓ�,�������E�"������=�Q�Jl��D���P�E�!�эU�R�E���C �u��E�P�E���C ���M�u��E���  �����������E�"�#�����=�Q�Jl��D���P�E�!�эU�R�E��C �E�P�E�    �E��yC ��=�E�    ���   ���   �E�P�E��у��E�    �$�����=�B�P`�M�Q�ҡ�=�H�Ad3�Wj��U�h0�R�Ћ�=�Q�J`�E�P�E�:�ы�=�B�PdWj��M�h$�Q�҃�(��=���   �Bx���E�;��P�M�Q������R�   �M�QP�������<R�]���  P�E�=耘 ��=�H�Al������R�]��Ћ�=�Q�Jl������P�E�;�ы�=�B�Pl�M�Q�E�:�ҡ�=�H�Al�U�R�E�0�Ѓ�,�������E�"裰����=�Q�Jl��D���P�E�!�эU�R�E��B �E�P�}��E���A ��=�}싑�   ���   �E�P�E��у��}�������=�H�A`�����R�Ћ�=�Q�Jdj j������h�P�э����R�E�>�q� ��=�H�Al�����R�E��Ѓ�3��� ���Q�� ��=���   ���   �M�Q�E��҃��������}��E��g= �������E� �X= �������E������F= �   �M�d�    Y_^[��]� ������������̡�=V�񋈜   ���   V�҃��    ^���������������V��V�@ ���    ^�������������U��Q3�9A~V�u�2@��;A|�^]� ���������������U��VW�}���}_3�^]� �F;ǋ���S�]��N�U��uh��hJ  �� ��[_3�^]� ��;��6  )^�F��   @����   h��+؋F��^�NÉF���u"��=�P�I���  ��hX  P�у��"��=�R���  �I�hY  �QP�҃��ȉ���j����F�@���F�N��~N+Ǎ@��R�U��+�@��P��@��P�u �E�N���+�R�@��RQ�}u ���  �U�@��P��+Í@��P�R��   ��~�V���Q�R�@��R�9u ���F��@���V�   �F�D������C��;^~k�h����u#��=�Q���  �[��hu  P�у��"��=�J�[�hv  �RP���  �Ѓ��ȉ���F����F�@���F�^�F;�}(�N+Ǎ@��R����E�R�@��P�wt ���} tF�N;�} ��+��@��R�I�N��j R�Js ���E�V�@��P���j P�+s ���} tP�N��;�}!�F�I����+х�t�P�P�����u�V����M��~��t�P�P�����u��؋E[�F_�   ^]� U��V��MW��|$�~;�}�> t�~ uh��h�  �� ��_3�^]� �E��;�|��蔚��_�   ^]� S�;�|�ߋ�+���;ȉ]��   ^��~�F�I��QP�[��P�/s ���N��~;ύI���V�  ������V+ӍR��R��)F+ȍ@�N�N�Q�+�Q��r �F��=�Q����  �@h���h�  �PQ�҃������   �N)^�I[��_�V�   ^]� �F+Ë^�D8�����W�@��;ʋ]�E}+�F+�+����R��R��R�I��R�Mr �E��;F}J��=�Q����  �@h���h�  �PQ�҃����u	[_3�^]� �N�I���E�F�V)^[_�   ^]� ���������U��S�]V���}^3�[]� �F;Ë���W�}�9�N�U��uh��hJ  �� ��_^3�[]� ��;��  )~�F��   @����   h��+��F��~�NǉF���u"��=�P��    ���  hX  P�у����=�R���  �hY  �QP�҃�����o����N�V���M�F��~>+���R��+�э�Rˍ�R��p �F�U��    Q+׍�QP��p ����   ��R��+׍�R��P��   ��~�V��    Q�R��R�p ���F����V�   �F�D������G��;~~f�h����u#��=�Q���  ��    hu  P�у��"��=�Jhv  ��    RP���  �Ѓ�����k����N���V�~�F;�} �N�U+���P��P���Q��o ���} t=�F;�}�N��+���R��j R�n ���E�V��    Q��j P�n ���M_�N^�   []� ���������������U��VW�}���|$�N;�}�> t�~ uh��h�  ��� ��_3�^]� �E��;�|���D���_�   ^]� S�;�|�ً�+���;��]��   ^��~�F��    QP��R��n ���N��~;ύ��V��   ������V+���R��)F+ȉN�N�Q�+�Q�n �F��=�Q����  h���h�  �PQ�҃������   �N)^[��_�V�   ^]� �F+ÍD���~�Q���C�^;�}!�U�F+�+���Q׍�Q��R�n ��;^}C��=�H����  h��h�  ��    RP�у����u	[_3�^]� �V���F�^�])^[_�   ^]� ��������������U�존=V��H�QV�ҋ�=�Q�M�R0QPV�҃���^]� ��������������U�존=�P�Ej PQ�J �у����@]� �������������U��Q�E;�u	�   ]� }+�RP����]� jj+�PR�.���]� ����������U��j�h!d�    P��V�'3�P�E�d�    �E�    ��=�H�A`�U�R�Ћ�=�Q�M�Rp�E�PQ�ҡ�=�H�A�U�R�E�   �Ћ�=�Q�MQ�J0P�E�P�ы�=�B�u�H`V�ы�=�B�Pp�M�VQ�ҡ�=�H�Al�U�R�E�   �E� �Ѓ�,�ƋM�d�    Y^��]��������U��V��W�~��}_3�^]� jjjW������t�F�M��_�   ^]� �������<���o �����U��V���<���o �Et	V�#a ����^]� ���������U��M�UV�uW��r�;u��������s��tE��9+�u1��v6�B�y+�u ��v%�B�y+�u��v�B�I+���_��^]�_3�^]�����������U��QV��j �M���Y �F���s@�F�M���Y ^��]�������U��QVW��j �M��Y �G��v	���sH�G�w����֍M�#��Y _��^��]�����H�����������U��QW�9��t=j �M��SY �G��v	���sH�GV�w����֍M�#��WY ��t
��j����^_��]����U���EV���H�t	V�_ ����^]� �������������̰�������������̸   �����������U��Q�A$V�0W�}j �M�E�    �7�X �F���s@�F�M�X ��_^��]� �U��j�hYd�    PQVW�'3�P�E�d�    ���E�    �u���E�    葽  ��=�H@�Q`VW�E�    �E�   �҃��ƋM�d�    Y_^��]� �����������̡�=�P�Bl��Q��Y��������������U��MV3���� ��t��=���   ���ȋB(�Ѕ�u��^]� ��������������U��j�h�d�    P��SVW�'3�P�E�d�    ���E�    �� �O ���EP�,h P���Ŀ �M�Q�������jh�  �M��E����  jh�  �M����  �URh�  �M����  jh�  �M���  ��=�H@�Adj�U�RV�Ћ]����3���� ��t��=���   ���ȋB(�Ѕ�u�WV���^� ��=���   �Bj j���ЍM��E� �{�  ��=�Q�Jl�EP�E������у��M�d�    Y_^[��]� �����������U��j�h�d�    P��4SVW�'3�P�E�d�    ��u�=�HT�U�A,j R�Ѓ��E��u�M�d�    Y_^[��]� �M�Q���� ���   +��   �]�ƨ   ���g������������E�    ;�r��n �N��i��   �T9Rh�  �M���  �N+N���g�����������;�r�n �N��9�    tIS���S  ��LPh�  �M��
�  �U���R�M��, �E�Ph�  �M��E���  �M��E� �Z, �M�Q�M�^� �M��E�������  �   �M�d�    Y_^[��]� ������U��j�h�d�    P��TSVW�'3�P�E�d�    ���}�=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�у����   +��   �]�Ǩ   ���g������������E�    ;�r�cm ��=�Q�R ��i��   Gj �M�Q��\P�ҋ�=�H�Al�ލU��R���E������Ѓ�����  ��=�QT�u�B,j	V��3Ƀ��E;�u3��M�d�    Y_^[��]� �M�M�h�  �M��E�   �n� j �M�QP���E��ܰ �M��E�耜 �E�   �E�    ��=���   �@�M�Q�U�R�E��Ћ�=���   �
�E�E�P�E��у��} tW�E�   �E�   h�  �M��E��� j �U�RP���E��p� �M��E���� ��=���   ��U�R�E��Ѓ��u�M�Q����� S���E�� Q  ��4Ph�  �M��?�  S���Q  ���    tIS����P  ��\Ph�  �M��U�  �U���R�M��f) �E�Ph�  �M��E��Q�  �M��E��) �M�Q���� �M��E��>�  ��=���   ��M�Q�E������҃��   �M�d�    Y_^[��]� �������U��j�hq�d�    P��TSVW�'3�P�E�d�    ���}�=�H�A`�U�R�Ћ�=�Q�Jd3�Sj��E�h��P�у����   +��   �u�Ǩ   ���g����������]�;�r�j ��=�Q�R ��i��   GS�M�Q��pP�ҋ�=�H�Al�ލU��R���E������Ѓ�;���  ��=�QT�u�B,jV�Ѓ��E;�u3��M�d�    Y_^[��]� �]�]�h�  �M��E�   褧 S�M�QP���E��� �M��E�跙 �E�   �]��=���   �@�M�Q�U�R�E��Ћ�=���   �
�؍E�P�E��у���tW�E�   �E�   �h�  �M؈]��� j �U�RP���E�譭 �M؈]��2� ��=���   ��U�R�E��Ѓ��]�M�Q���:� �uV���E��[N  ���    tIV���JN  ��pPh�  �M�詼  �U���R�M��& �E�Ph�  �M��E�襼  �M��E���& �M�Q����� �M��E�蒵  ��=���   ��M�Q�E������҃��   �M�d�    Y_^[��]� �����������U��j�h܀d�    P��TSVW�'3�P�E�d�    ���}�=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�у����   +��   �]�Ǩ   ���g������������E�    ;�r��g ��=�Q�R ��i��   Gj �M�Q��pP�ҋ�=�H�Al�ލU��R���E������Ѓ����  ��=�QT�u�B,jV��3Ƀ��E;�u3��M�d�    Y_^[��]� �M�M�h�  �M��E�   �� j �M�QP���E��\� �M��E�� � �E�   �E�    ��=���   �@�M�Q�U�R�E��Ћ�=���   �
�E�E�P�E��у��} tW�E�   �E�   h�  �M��E��b� j �U�RP���E��� �M��E��t� ��=���   ��U�R�E��Ѓ��M�Q�M�~� S���K  �@l�5���E�   �]�E�]�h  �M��E��� j �U�RP���E��z� �M��E���� ��=���   ��U�R�E��Ѓ�S���<K  ���    tIS���+K  ��pPh�  �M�芹  �M���Q�M��# �U�Rh�  �M��E�	膹  �M��E���# �M�E�P��� �M��E��r�  ��=���   �
�E�P�E������у��   �M�d�    Y_^[��]� �����������U��j�hG�d�    P��TSVW�'3�P�E�d�    ���}衴=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�у����   +��   �u�Ǩ   ���g������������E�    ;�r��d ��=�Q�R ��i��   Gj �M�Q��P�ҋ�=�H�Al�ލU��R���E������Ѓ��   ����  ��=�QT�u�B,jV��3Ƀ��E;�u3��M�d�    Y_^[��]� �M��M�h�  �M؉]��͡ j �M�QP���E��;� �M؈]���� �E�   �E�    ��=���   �@�M�Q�U�R�E��Ћ�=���   �
�E��E�P�]��у��}� tR�E�   �]�h�  �M��E��G� j �U�RP���E��է �M��E��Y� ��=���   ��U�R�]��Ѓ��M�Q�M�d� �E�   �]�h�  �M��E��� j �U�RP���E��w� �M��E���� ��=���   ��U�R�E��Ћu��V���6H  ���    tIV���%H  ��Ph�  �M�脶  �M��Q�M��  �U�Rh�  �M��E�	耶  �M��E���  �M�E�P��� �M��]��m�  ��=���   �
�E�P�E������у��ËM�d�    Y_^[��]� ���������U��j�hЁd�    P���  �'3ŉE�SVWP�E�d�    ����j ��ٕH�����T���ٕL�����H�����PٝP��������Q�����ٕ���R�荅8���ٕ���3�ٝ���P��������X���ٕ ���ٕ���ٕ���ٕ8���ٕ<���ٝ@���������=�Q�J`��4���P�ы�=�B�PdVj���4���hp�Q�ҍ�4���P�u��z ��=�Q�Jl��4���P�E������ы��   +��   �����������������\�����
  ��`������   +��   ���������������9�\���r��` ���   �`����{ �   ��x������   ��=�B�P`��4���Q�ҡ�=�H�Idj j���x���R��4���P�у���T�����4���R�E�   �TX ��D�����=�H�Al��4���R�E������Ѓ���D��� t��D���Q�k� ���U܋E�RP�� ������h�������	  ���   +��   ���������������9�\���r��_ ��=�B���   �P`�`��������Q�ҡ�=�H�Adj j������WR�Ѓ���=���   �R|�����P���E�   �ҡ�=�H�Al�����R�E������Ћ�=�QH�B|j h�  V�Ћ�=�QHj ��t����B|h�  V�Ѓ��}� ǅp���    ~o3��
��$    �I �U�t��X���+���d����t+���l����t�+׉��l���+��p�P��d����P��p���B�� ��;U܉�p���|���h���3�9}���   ��X���م����م������t���م�����Rم�����م����ҋ��   م������G��؅�������@؍���������H��ٝt���م�����؅�����@�������H��ٝl���م�����؅�����@�������H��ٝd���مt���ٝH�����H���مl����A�ٝL�����L���مd����A�ٝP�����P����A�;}��>������������؃; ��  �}� ��  ��M�ٕ����Qٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٕ����ٝ�����1� ������l������"  �}� ǅd���    �  3���p������p����M�T�t�|���   �<�<���t�����p����L�I�R���4v�4������P����H�@��T�����X�����t������\����H�@��`������h����N��d����F��p����J��l�����R��x�����t�����|����   ��P���������󥋍l���葩 ��=�QD��d����RX������QVP�҃�p��� F��;u܉�d����������l�����h���j W��蔱 ��=���   �Bj j����j h�  ��� � ����   ��=�Q�J`�����P�ы�=�B�Pd3�Wj������hH�Q�҃���=���   �Bx���E�   ��P�����Q�����R����P�E��:s ��=�H�Al�����R�E��Ћ�=�Q�Jl�����P�E������у��3�9{��  ��=�B�P`��$���Q�ҡ�=�H�AdWj���$���h��R�Ѓ����   +��   ���g����������ʃ����   �E�   ���g�un+��   ��$���R����������u�Z ���   ��=�B����t����H`����l���W�ы�=�B��t����PpWQ�҃�V��������  +��   ������������  ��$���Q���   +��   ���g�����������u��Y ���   ��=�B����t����H`����l���W�ы�=�B��t����PpWQ�҃�V���������   +��   ���g�����������   �;��?  ǅp����   h)  �� ��=�Q������l������/  �J`��@���P�ы�=�B�Pdj j���@���h<�Q�ҍ� ���WP�E��6� P��@���Q��0���R�E��>�����=�Q�Rp��$���QP�E��ҡ�=�H�Al��0���R�E��Ћ�=�Q�Jl�� ���P�E��ы�=�B�Pl��@���Q�E��ҡ�=���   �R|��<��$���P���ҋ��� 3�9u܉�t���~�E�9<�u��t���V�� F;u�|拍h���3��C� ��t��=���   ���ȋB(�Ѕ�u狍h���V��l���V賭 ��=���   �Bj j���Ѝ�$���Q���   +��   ���g�����������;�r��W ��=�Q���   �p������ĉ�t�����t���P�B`�Ћ�=��t����Q�JpPV�ы�h�����R����������   +��   ��p����   ���g����������G�;��������h���3���=�Q�Jl��$���P�E������у���T���WWWV��K ��=���   �PWj���҉������������������������� ���ǅ����   ��������T���������Qh�   �E�	   ��������������o ���E���������������   �U��X���订  ���   +��   ��\�����`���x��������������F�\���;��@����   �M�d�    Y_^[�M�3���I ��]ËJl��$���P�E������у�3����3�  3������������������U��j�h �d�    P��SVW�'3�P�E�d�    �񋎸   +��   ���g����������3���-  �]����   +��   ���g�����������;�r�{U ���   E��N P�2M ����uihG  �R� ��������   ���   +��   ���g�����������;�r�$U ��=���   ���   E��R|P���ҋN j j W�I WS������WS��������~ W��Su�b��������WS���r���jj���� ��=���   �Bj j���Ћ��   +��   �E�   ���g����������C�;�������   �M�d�    Y_^[��]Ë�=�B�P`�M�Q�ҡ�=�H�Adj j��U�h��R�ЍM�Q�E�    ��k ��=�B�Pl�M�Q�E������҃�3��M�d�    Y_^[��]����������������U��j�hR�d�    PQSV�'3�P�E�d�    ��u����   P�E�   �A ���   P�A �����   ��y  ���   3�;�t	P�'A �����   P���   ���   ���   �A ���N\�E��w �N@�E��k �N$�]��` ��=�H�Ql��V�E������҃��M�d�    Y^[��]�����U��j�h��d�    P��SVW�'3�P�E�d�    ��u��=�Q�FP�B`�Ѓ��N$�E�    �/ �N@�E��# �N\�E�� ���   ���E�薃  ���   ���E�腃  3��Fx�F|���   ǆ�   �����G�E��E�9Gv�PR ��M��O�M�;Ov�;R �M��U�R�U�RQP�E�P���jb  �{9{v�R ��M��K�M�;Kv��Q �M�U��WRQP�E�P����o  �ƋM�d�    Y_^[��]��������������U��j�h�d�    P��\  �'3ŉE�SVWP�E�d�    �u�ٿ   W��0���謌  j@WV��8����E�    超  ��u+��0����H��8�����0������y( u��j P�gu  ������ ��  ��=�Q�J`������P�ы�=�B�Pdj j�������h��Q�ҡ�=�H�A`������R�E��Ћ�=�Q�Jdj j�������h �P�ы�=�B�P`������Q�E��ҡ�=�H�Adj j�������VR�Ѝ�����Q������R������P�]�������H������QP�� ���R�E�����P�E��+h ��=�H�Al�� ���R�E��Ћ�=�]��Q�Jl�����P�ы�=�B�Pl������Q�E��ҡ�=�H�Al������R�E��Ћ�=�Q�Jl������P�E� �у�$�������E������,�  ������Rǅ����P���: ��3��F  ��=�H�A`������R�Ћ�=�Q�Jdj j�������h��P�э�����R�E��
h ��=�H�Al������R�E� �Ћ�0����A��8��������c  j
��0����xv  ��Rjc������P��0�����  j������Qh<���Z ����uG{|���   +��   ���   ���������������;�r�N ���   ����+΍D�h��  j������Ph���mZ ����uJ��   ���   +��   ���   ���������������;�r�XN ���   ����+֍D�l�_  j������Qh���	Z �����  ��   ���   jx������@j R�������:E ��l���   ������󥋍�������   Q����  ���   +��   ���   ���������������;�r�M ���   ����+�3��|�d���   +��   ���   ���������������;�r�lM ���   ����+Ή|�h���   +��   ���   ���������������;�r�-M ���   ����+Ή|�l�   �4j������Ph����X ����u���   {xQ���   ��1  ��d8��0����B��8����������8����k  ��u+��0����H��8�����0������y( u��j P�p  �s|3ɋƺ   �������Q�9 �����t�V���|�H�Q�����Q��Q�y��3����   �؉��   3ɋƺ   �������Q��8 ����t!�V���|��H�Q�����Q��Q�y����3����   ���   +��   ��������������3���C  3����   +��   ���������������;�r�K ���   ǋ@d3�@�    �������Q�-8 ���   +��   ���������������������;�r�SK ���   �������Tp���   +��   ���������������;�r�K ���   ǋ@d3�@�   �������Q�7 ���   +��   ���������������������;�r��J ���   �������T9t���   +��   ��������������F�x;�������������E�������{  ������Qǅ����P��|5 ���   �M�d�    Y_^[�M�3���= ��]� ��������U��j�hÄd�    P��l  �'3ŉE�SVWP�E�d�    ��j�������#�  �������^\P���E�    �� ��=�Q�JP������jP�E��ы�=���B��H  hȩGh�  W�ы�=�JjWP�������������ATR�Ћ�������$j@jQ�������}  ��u+�������J���������������y( u��j P�jm  ������ ��  ��=�H�A`��p���R�Ћ�=�Q�Jdj j���p���h��P�ы�=�B�P`��`���Q�E��ҡ�=�H�Adj j���`���h �R�Ѓ�(��(���Q���E�� P��`���R�� ���P�E��������p���QP������R�]�����P�E��U` ��=�H�Al�����R�]��Ћ�=�Q�Jl�� ���P�E��ы�=�B�Pl��(���Q�E��ҡ�=�H�Al��`���R�E��Ћ�=�Q�Jl��p���P�E��ы�=�B�Pl������Q�E� �҃�4�� ����E������=y  �� ���Pǅ ���P���2 ��3��r  ��=�Q�J`��`���P�ы�=�B�Pdj j���`���h��Q�ҡ�=�H�A`��p���R�E��Ћ�=�Q�Jdj j���p���h �P�у�(�����R���E��/ P��p���P�� ���Q�E�	�W�����`���RP��(���P�E�
�?���P�E���^ ��=�Q�Jl��(���P�E�
�ы�=�B�Pl�� ���Q�E�	�ҡ�=�H�Al�����R�E����E���=�Q�Jl��p���P�ы�=�B�Pl��`���Q�E��ҋ������@��������0�������  �l�������������$    �d$ ������j
�������m  ��Qh�   ������R�������!�  j������Ph���Q �����  ��   �Ô   ��G��������������+  �O���   Q����x  ������R������h��P��R ��=�Q�J`��p���P�ы�=�B�@dj j�������Q��p���R�Ѓ� �K+K���g������������E�;�r�SE �C�������=�JP�Ap��p���R�Ћ�=�Q�Jl��p���P�E��ыK+K���g�����������;�r��D �K������Ǆ
�       ��  j������Ph���P ����������u^�����Qh��R��Q ���   +��   ���g�����������;�r�D ݅������   ٝ����م�����\�q  jRh���,P ����ud�����P������h��Q�gQ ���   +��   ���g�����������;�r�D ݅������   ٝ����م�����\��  j������Rh���O ����u)W���   ��(  ��P������h��P��P ���  j������Qh���kO ������   ��X���R��H���P��P���Q������hp�R�P ݅P�����ٝ�������   W���|(  م�����XW݅H�����ٝ�����_(  م����W�X ��݅X���ٝ�����B(  م�����X$�  j������Phl���N ������   ��X���Q��H���R��P���P������h\�Q��O ݅P�����ٝ�������   W����'  م�����X(W݅H�����ٝ�����'  م����W�X,��݅X���ٝ�����'  م�����X0�d  j������RhX��N ������   ��X���P��H���Q��P���R������hH�P�BO ݅P�����ٝ�������   W���*'  م�����X4W݅H�����ٝ�����'  م����W�X8��݅X���ٝ������&  م�����X<�  j������QhD��pM ������   ��X���R��H���P��P���Q������h4�R�N ݅P�����ٝ�������   W���&  م�����X@W݅H�����ٝ�����d&  م����W�XD��݅X���ٝ�����G&  م�����XH�  j������Ph,���L ����uZ������Q������h �R�N ��j ������P������� N��������Q���   W���E���%  �ȃ�L�]`���������vj������Ph��SL ������   ������Q������h�R�M ��j ������P�������M��������Q���   W���E��_%  �ȃ�\��_����������=�B�PlQ�E��҃�W���1%  ǀ�      �������@�������������������^  ��u+�������I���������������y( u��j P��c  j��D����z  ��4����^@R���E��t�  ��=�H�AP��4���jR�E��Ћ�=�Q����H  hȩGh7  W�Ћ�=�Q�JTjWP��������4���P�ы�������$j@jR��L����Ss  ��u+��D����H��L�����D������y( u��j P�c  ������ ��=�Q�J`��`���P��  �ы�=�B�Pdj j���`���h��Q�ҡ�=�H�A`��p���R�E��Ћ�=�Q�Jdj j���p���h �P�у�(�����R���E��I�  P��p���P�� ���Q�E��q�����`���RP��(����P�]��X���P�E���U ��=�Q�Jl��(���P�]��ы�=�B�Pl�� ���Q�E��ҡ�=�H�Al�����R�E��Ћ�=�Q��p����E�P�Jl�ы�=�B�Pl��`���Q�E��ҡ�=�H�Al��4���R�E��Ѓ�4�������E���n  �������P�Q�������p( ��=�B�Pl������Q�E� �҃��� ����E������n  �� ���P�� ����0( ��3���  �ы�=�B�Pdj j���`���h��Q�ҡ�=�H�A`��p���R�E��Ћ�=�Q�Jdj j���p���h �P�у�(�����R���E���  P��p���P�� ���Q�E��������`���RP��(����P�]�����P�E��BT ��=�Q�Jl��(���P�]��ы�=�B�Pl�� ���Q�E��ҡ�=�H�Al�����R�E��Ћ�=�Q��p����E�P�Jl�ы�=�B�Pl��`���Q�E��ҋ�D����@3���0��L�����������  j
��D����c  ��Qh�   ������R��D����x  ���   +��   ���g����������3����   ��������=�Q�J`��p���P�ы�=�B�@dj j�������Q��p���R�Ѓ����   +��   ���g������������E�;�r�; ��=�J���   �����j ��p���RP�A �Ћ�=�Q�Jl���ߍ�p����PG�E��у���u4���   +��   �������   ���g����������C�;������������������j������Qh���NF �����*  ���   +��   ���g�����������;�r�A: ���   i��   �TlR������h�P�SG ��D����I��j
��D����^a  ��Rh�   ������P��D�����v  ��=�Q�J`��`���P�ы�=�B�@dj j�������Q��`���R�Ѓ����   +��   ���g������������E�9�����r�9 ���   ��=�H�Ap�|p��`���WR�Ћ�=�Q�Jl��`���P�E��ы�������   j	������Rh��E ������   ��D����Hj
��D����c`  ��Qh�   ������R��D�����u  ��=�H�A`��8���R�Ћ�=�Q�Rdj j�������P��8���Q�҃����   +��   ���g������������E�;�r�8 ���   ��iɔ   ���   ��=�Q�JpP��8���P�ы�=�B�Pl��8���Q�E��҃���D����@��L����b���3���L���9�����t ����H  ��u3�������Q�cC ����t3���T�����\�����X�����d�����h�����`�����l�����p�����=��t�����x���ƅ���� ƅ���� ��|�����������X�����h�����x�����T�����d�����t���������������������;�u)��D����H��L�����D�����9y(u��WP�f[  ������V��C ������Y  ��=�Q�J`������P�ы�=�B�PdWj�������h̨Q�ҡ�=�H�A`������R�E��Ћ�=�Q�JdWj�������h �P�ы�=�B�P`��8���Q�E��ҡ�=�H�AdWj���8���VR�Ѝ�8���Q������R������P�E� ������H������QP�������!R�]�����P�E�"�"N ��=�H�Al������R�]��Ћ�=�E� �Q�Jl������P�ы�=�B�Pl��8���Q�E��ҡ�=�H�Al������R�E��Ћ�=�Q�Jl������P�E��у�$��=�B�Pl��4���Q�E��҃��������E��
g  �������P�P�������  ��=�Q�Jl������P�E� �у��� ����E�������f  �� ���R�� ����a  ���   �M�d�    Y_^[�M�3��( ��]����������������V��������������   ^�����������U��j�h�d�    P��$SVW�'3�P�E�d�    3��u�M�u���e  �E�]jV�M�Q�ˉu��E�   �E��*  �������   �U�U��    ��+�PV�M�Q���L  �MP�E�   �{  �}��E� r�U�R��! ��j�wV�EP���)  �����u�PV�M�Q���dL  �uP���E�   �B{  �}�r�U�R�! ���ƋM�d�    Y_^[��]� �E�M�d�    Y_^[��]� ���U��j�hM�d�    P��  �'3ŉE�SVWP�E�d�    �]����������������@����d  3��������u��d  j�������E��n  j@jS�������E��g  ��u)�������H��������������9q(u��VP�TW  9�������  ��=�Q�J`��d���P�ы�=�B�PdVj���d���h��Q�ҡ�=�H�A`��T���R�E��Ћ�=�Q�JdVj���T���h �P�ы�=�B�P`������Q�E��ҡ�=�H�AdVj�������SR�Ѝ�����Q��T���R��(���P�E�袽����H��d���QP��D����R�]�膽��P�E��J ��=�H�Al��D���R�]��Ћ�=�E��Q�Jl��(���P�ы�=�B�Pl������Q�E��ҡ�=�H�Al��T���R�E��Ћ�=�Q�Jl��d���P�E��у�$�������E�� c  ������Rǅ����P�� ���������|h  �������qh  3��  ��=�H�A`��d���R�Ћ�=�Q�JdVj���d���h��P�ы�=�B�P`��T���Q�E��ҡ�=�H�AdVj���T���ht�R�Ћ�=�Q�J`������P�E�	�ы�=�B�PdVj�������SQ�ҍ�����P��T���Q��(���R�E�
������H��d���QP��D����R�]�����P�E��~H ��=�H�Al��D���R�]��Ћ�=�E�
�Q�Jl��(���P�ы�=�B�Pl������Q�E�	�ҡ�=�H�Al��T���R�E��Ћ�=�Q�Jl��d���P�E��ы�=�B�P`��l������Q�������������ҡ�=�H�A`������R�E��������Ћ�=�Q�JdVS������hd�P�э�����R�E��fH ��=�H�Al��������@R�E��Ћ������A������������	  3ۉ������������j
��������V  ��Rh�   ������P�������Wl  j������Qh���; ������   ������R������hX�P�L< ��@�����Q��t�����  ��t����w\R���E���  ��t����E���  ���Q�  ������P��t����_�  ��t���Q���E���  ��t����E����  ��  j������Rh���g: ������  ��=�H�A`������R�Ѓ��������������E���;�v�P. ��������������������;�v�3. ������SVWQ��\���R�������@g  �   3�������������������ƅx��� �P�@��u�+�P������P��t����9  jj��t���Q��l����E���i  �   9�����r��x���R�N ��������P�� �ĉ8�p�x������������ƅx��� �������@ �� ��l����̉�����R�E��/s  ������P�E���u  ������������+θ�$I����������ʃ�H��w�- ������9^4r�v ��� ��=�B�P`��D���Q�ҡ�=�H�AdWj���D���VR�Ћ�=�Q�Rp������P��D���Q�E��ҡ�=�H�Al��D���R�E��Ћ��������   +��   �ƨ   ���g������������ �tw3ۍ�$    �N+N���g�����������;�r�E, ��=�Q�F�R j �������QP�҃����   �N+N���g����������GÔ   ;�r��N+N���g������������   �|
�̉�������  W����^  �N+N���g���ыN+N������x����g�����������;�r�+ ��=i��   ~�Q�Jp������WP�ыN+N���g�����������L��������������E��'  ������Rǅ����P��4 ��=�H�Al������R�E��Ѓ��*  �������j������Qh���6 ����u9������@P���   �������������  P������hP�R��7 ����  j������Ph<��i6 ������   ��0���Q��|���R������P������h@�Q�7 ݅����������ٝ�������   م��������   ݅|�����ٝ������م�����\����   ݅0���ٝ����م�����������\��/  j������Ph���5 ������   ��8���Q�� ���R������h4�P��6 ��l���Q��8���R�� ���P������h$�Q��6 ݅ ������   ٝ����م������$����   ���ܥ8���ٝ����م�����\����   ݅l���ٝ����م�����������\��f  j������Rh����4 �����H  ���������t������P���   ��  �Ht���������������c  ������P��P�����@  jj��P���Q��l����E���d  ��P�����-  ������R�� �ĉ0�@   �p�������@ �� ��l����̉�����P�E��>n  ������Q�E��q  ��H������� c  ��������������+˸�$I�����������   �;��L  �����������   ��������$    ������j/V�������\  P��x���R�������P�������E��h  ��x����E��^  j �������!  �xr�@���P��4 �X����������ǐ   P���s  �Hp�������\�j��������  �Hj h��Qj ���  ��tJj�������  �xr�@���P�}4 ��������R�ύX��  �������@p���Ή\���������������������+˸�$I����������F�;������+���$I�������������   j �������  �xr�@���P��3 ���������������������ǐ   Q�ύX����\  �Pph��j�������\2��  P�,  ����t<j�������  �xr�@���P�r3 �X���������P���  �Hp�\1�������������E��E"  ������Rǅ����P��� ��������������3��������@�������7���������9�����t ���r6  ��u3�������Q��0 ����t3���������������������������������������������������=������������ƅ���� ƅ���� ������������������������������������������������������������������;�u)�������H��������������9q(u��VP��H  ��=�Q�Jl��l���P�E��у��������E���U  ������Rǅ����P�� ��������;�t*������Q������������RQP�?G  ������R�� ��������P�������������������� ��������;�t*������Q������������RQP��F  ������R� ��������P�������������������} ���   �M�d�    Y_^[�M�3��I ��]� �������U��j�h��d�    P��<  �'3ŉE�SVWP�E�d�    �}�E��j j	�ωF ��r  j j�ω�r  j j�ωF�r  j j
�ωF��r  �F��=�Q�J`������P�у�������Rj������P���E�    ��s  ��=�R�NQP�Bp�E��Ћ�=�Q�Jl������P�E� �ы�=�B�Pl������Q�E������ҡ�=�H�A`������R�Ѓ�������Qj������R���E�   �is  �E�P�������9�  �������^$P���E��4�  �������E��u�  ��=�Q�Jl������P�E��ы�=�B�Pl������Q�E������҃�h����������  ������P���E�   ���  �������E�������  ��=�Q�J`������P�у�������Rj������P���E�   �r  P�������E��`�  �������~@Q���E��[�  �������E���  ��=�B�Pl������Q�E��ҡ�=�H�E������Al������R�Ѓ�h�����������  ������Q���E�	   ��  ����������}��/�  j�������"\  ������R���E�
   ���  ��=�Q�RTj h�   ������QP�E��ҡ�=�H�Al������R�E�
�Ѓ�j@j������Q��������T  ��u+�������J���������������y( u��j P�D  ����� ��=�H�A`�V  ������R�Ћ�=�Q�Jdj W������h��P�ы�=�B�P`������Q�E��ҡ�=�H�Adj W������h �R�Ѓ�(������Q���E����  P������R������P�E������������QP��d����R�]�����P�E��y7 ��=�H�Al��d���R�]��Ћ�=�Q�Jl������P�E��ы�=�B�Pl������Q�E��ҡ�=�H�E��Al������R�Ћ�=�Q�Jl������P�E�
�у�0������}��~P  �����Rǅ���P��
 ��3��  ������R�Ћ�=�Q�Jdj W������h��P�ы�=�B�P`������Q�E��ҡ�=�H�Adj W������ht�R�Ѓ�(��d���Q���E��~�  P������R������P�E�覩��������QP�������R�]�荩��P�E��#6 ��=�H�Al������R�]��Ћ�=�Q�Jl������P�E��ы�=�B�Pl��d���Q�E��ҡ�=�H�E��Al������R�Ћ�=�Q�Jl������P�E�
�ы������J��0j
�������E  ��Ph�   ������Q�������Z  �������<  ��u+�������J���������������y( u��j P�A  ������P��) ��;��`  ��=�Q�J`������P�ы�=�B�Pdj W������h̨Q�ҡ�=�H�A`��t���R�E��Ћ�=�Q�Jdj W��t���h �P�ы�=�B�P`������Q�E��ҡ�=�H�Idj W������R������P�э�����R��t���P��T���Q�E��ǧ����H������RP��D����P�]�諧��P�E��A4 ��=�Q�Jl��D���P�]����E���=�B�Pl��T���Q�ҡ�=�H�Al������R�E��Ћ�=�Q�Jl��t���P�E��ы�=�B�Pl������Q�E�
�҃�$�^4 ������P������������Q��������~ t/���   +��   ���g�����������t���d������������6�����3 j h  �4 ��������}���L  �����Qǅ���P��l ���   �M�d�    Y_^[�M�3��� ��]� ��������Q�P��2 Y��̋A��P�D
�X���U��V��N+N��������������W�}�;�r�� �V����+�_��^]� �U��V��N+N���g����������W�}�;�r� ��i��   F_^]� ���U��V��N+N��$I����������W�}�;�r�[ �V��    +�_��^]� ���������������U��V���ŧ���Et	V�� ����^]� ���������������U��j�h��d�    PQV�'3�P�E�d�    ��u�=�H�Q`V�����V$�FL�V P�V�E�    �V0�V,�V(�V<�V8�V4�VH�VD�^@��=�Q�B`�Ћ�=�Q�F\P�B`�E��Ћ�=�Q�FpP�B`�E��Ћ�=�Q�J`���   P�E��у��ƋM�d�    Y^��]�U��j�h��d�    PQV�'3�P�E�d�    ��u�=�H�Al���   R�E�   �Ћ�=�Q�Jl�FpP�E��ы�=�B�Pl�N\Q�E��ҡ�=�H�Al�VLR�E� �Ћ�=�Q�BlV�E������Ѓ��M�d�    Y^��]���U��V��V�P�� ���Et	V� ����^]� �����U��A�U��Q �E��U+ЋA0�]� ��������������̋A �8 t�I0��3�����������������U��A�U��Q$�E��U+ЋA4�]� ���������������V���F@t�F�Q�l ���V�    �F �     �N0�    �V�    �F$�     �N4�    �f@��F<    ^�������U��Q�A8V�0W�}j �M�E�    �7�W� �F���s@�F�M�k� ��_^��]� ̍Q�Q �Q�Q$�A�A�Q(�Q0�A�A�Q,�Q4�     �A$�     �Q4�    �A�     �Q �    �A0�     ���������U��j�hI�d�    PQSVW�'3�P�E�d�    ��u�=�H�Q`V�ҡ�=�H�}�QpVW���G�^�^L�GS�^�G�F�O�N�W �V �G$�F$�O(�N(�W,�V,�G0�F0�O4�N4�W8�V8�G<�F<�O@�N@�WD�VD�GH�FH��=�Q�B`�E�    �Ћ�=�Q�Jp�GLSP�ы�=�B�H`�^\S�E��ы�=�B�Pp�O\SQ���Gl�^l��=�H�Q`�^p�E�S�ҡ�=�H�Ap�WpSR�Ћ�=�Q�B`���   S�E��Ћ�=�Q�Jp���   SP�ы��   ��<���   �ƋM�d�    Y_^[��]� �����U��VW�����u�E ���t��3ҋE����+��G����;Bw��t�	�3�;As� w��_^]� ���������U��VW�����u�� ���t��3ҋE�4�    +��G���;Bw��t�	�3�;As� w��_^]� ���������U��M����w3ɋ���+����R�  ����]Ã��3����xsڍEP�M��E    �� h���M�Q�E�<��J ���U��M����w3�iɔ   Q���  ����]Ã��3���=�   sߍEP�M��E    � h���M�Q�E�<��� ��������U��M����w3ɍ�    +���R�^�  ����]Ã��3����sڍEP�M��E    �> h���M�Q�E�<�� ���U��EVP���j �<���^]� ����U�존=VW�}��H�QpVW���G�^�G�^�G�F�O�N�W �V �G$�F$�O(�N(�W,�V,�G0�F0�O4�N4�W8�V8�G<�F<�O@�N@�WD�VD�GH�FH��=�Q�Rp�FLP�OLQ�ҡ�=�H�Ip�V\R�G\P���Gl�^l��=�B�@p�NpQ�WpR�Ћ�=�Q�Rp���   P���   Q�ҋ��   ��(���   _��^]� ���U��S�]V�u;�t#W�}V��������Ɣ   �ǔ   ;�u��_^[]ËE^[]��������U��S�]V�u;�t#W�}��   ��   V������;�u��_^[]ËE^[]��������U��E��V��M�Q�F�h��� ��V�H�N�P�V�@�F����^��]� ���������������U���E��QP��� ��]� ��������U��S�]V�u;�tW�y�WP�� �F��;�u�_��^[]� U���E��QP��� ��]� ��������U��S�]V�u;�tW�y�WP�� �F��;�u�_��^[]� U��E]� ������U��E�UV�1W��+�W�}WP�FR��_^]� �������������U��S�]VW�}��+�9us� �E�MVSPQ� ����_^[]� �����������U��E]� ������U��E�UV�1W��+�W�}W�}WP�F(R��_^]� ���������U��S�]VW�}��+�9us� �E�MVSPQ� ����_^[]� �����������U��V��F�h���~�FP�7 �}�NQ��  ���E�H�t	V�b�  ����^]� �������̋��Q�D(��t�H�� ���������V��W�~8�����t������W��  ��_�N^��� ����̃��� ���������̃���������������U��U��@R�Uj�R��]� �������̋�� �����������3���������������� ������������̋A$�8 t�I4��3�����������������V���P�҃��u�^ËF0��F ��Q��^����������U��E����3ɉH�H�H]� ���U��E����3ɉH�H�H]�  ���U��A � ��t<�Q;v5�U���t:P�t�A@u"�A0� �A ����t�A ����]� 3�]� ���]� ̋Q V�2��u���^�SW�y0����;�s�_[^��A@u/�A$� ��t&;�w9q<v9A<s�A<��A<+�I ��_[^�_[���^����������������U��SV�q$�W��t9A<s�A<�]����   �A �����   �E��u�A�y<+8�u��'��u��u�A�u��+8����t�5����u����   �A� �y<+�;���   +Q0�)�Q ����   �Q$�����   �Q4�ЋA R��AR�R������p��te���t_�E�=����u�A�Y<+�u����u�A�u��+��	����u�u��|�A� �Y<+�;�+Q4�)�I$�
����5���E_3ɉ0^�H�H�H[]� ��U��E�UVW�y$�4���t9A<s�A<���;���   S�]$��tR�Q ���tI��|w�A� �y<+�;�d+Q0�)�Q ��tX�Q$���tO�Q4�ЋA R��AR�R�����4��t-�?��t'��|#�A� �Q<+�;��Q4+��)�I$������[�E3�_�0�H�H�H^]�  ��������������U��V�q���Q�F�D�X�P� P��[� ���Et	V���  ����^]� ����U��V��W�~8�����t��襘��W��  ���N�h� �Et	V��  ��_��^]� �������������U��V��W��������~8�����t���J���W�T�  ���N�� �Et	V�=�  ��_��^]� ��U��Q�U�E�M���u	;A��   SVW�y;�st+�;�wn�   +���yr
���M�	����M��E�WQS�� ������t5�U�ERPV诖������t,�M�+ލ|�WR�^S� ������u�_^���[��]� �E��x�Mr�	_��^+�[��]� �U��SV�uW��9ws��� �G+Ƌu;�s���]��;�r�Ãr�����MP�EP�W��������u;�s
_^���[]� 3�;���_^[]� �U��M����w3�Q���  ����]� ���3����s�EP�M��E    �� h���M�Q�E�<��	 ��������������V�����t(��u�� ��xr�H��H�@�9Fr�� �F^����������U��E��u&�yr�I�E�U�]� �E�U���]� �yr�I����UP�EP�Q�� ��]� ���������U��j�h{�d�    P��SVW�'3�P�E�d�    �ى]�K����o� j�E�    ��  ������t.�� ���� j �M������ �G���s@�G�M��� �3��ˉs8�����ËM�d�    Y_^[��]�U��S�]V�uW���    ��t)��t%�V�F��r����;�w��r� �N�;�v�q �7�_��_^[]� ������������U��E�M�UV�uPQRV�N ����^]����������������U��E�M�U ��E��   ]� ����U��E�M��   ]� ������������U��E+E�M;�s��]� ����������U��S�]V�u��+θ����������������+ȋE�ȉM��;�t#+�W��I �<���x�   �;�u�E_^[]�^��[]����������������U��S�]V�u��+˸����������������+���ɋыM��+�;�t+�W�M��M��x�<�   ���;�u�_^[]����������������U����US�]V�uW�}2��E��M��E��E�PQRWVS����+��g�����������iɔ   ����_^+�[��]��������U��U�ES�];�tVW��t�   �����x��x;�u�_^[]����������������V��F � ��t=�N0�	��~�F0��F � �V �� ^Å�t�N0�9 ~����F ��Q���	��P���҃��u�^ËF �8 t�N0�9 ~��^Ë�P��^������U��QV3�9uW���u�~nS�]��������~6�M;ȋ�}��G ��UVQRS� �G0)0u�)u�G ރ�0�u����P���҃��tF�C�M�u��} �[_��^��]� _��^��]� ������U��QV3�9uW���u�~mS�]���3�����~3�M;ȋ�}��VSP�G$�Q� �G4)0u�)u�G$ރ�0�u����P�B���Ѓ��tFC�M�u��} �[_��^��]� _��^��]� �������U��j�h��d�    PQVW�'3�P�E�d�    �M��A��P�D
����q����E�    �������~8�����t���ߐ��W���  ���N�� �F��H�D1�X��M�d�    Y_^��]����������������U���V���F@Wt �~$���t�N<;�s�F4� +��N4��E���u
_3�^��]� �V$�:S��t$�N4����;�s�	�v$�[�Q�_�^��]� �F@u=��u3���F4�N�+ߋ���� s�    ���v������+�;�s��u��u[_���^��]� �P�ND�E���������F��M���vSQ�M�QW������M�����u"�V�~<�:�F$�8�V4�E���F@u7�GPW�V�F$��+�V<� �V��+�+��V$ǉ��+�U��F4��F@t�V�:�F �     �V0�:��F$��F BR�+��RW���?����M��F@t	Q�0�  ���F4�N@��v$��A��E[_�^��]� �����������̋P���  Y�������U��S�]V��W9^s�a� �F�}+�;�s����v^�N��r�V��V�U��r�V��V+�P�E��P+�Q�R�0� �F+ǃ��~�Fr�N_� ��^[]� �N� _��^[]� ��U��} VW�}��t'�~r!�FS���vWSjP�� ��S�-�  ��[�~�F   �D> _^]� ����U��E�MPQ�D 3҃������]�V��~L t#��Pj��҃��t�FLP� ����}���^�3�^�U��A � S�]��t,�Q9s%���t�@�;�u�A0� �I �	��@���#�[]� �AL��t$���t�y< u��PQ� �����t��[]� ���[]� �V��F ���t�Ћ�V0��;�s�^Ë�PW���ҋ����u_�^Ë�PW���ҋ�_^������������U��V��NLW��tl�U�}��u	��u�G�3�WPRQ�n ����uG�~L���FH�FA�������t�G�F�F�G�~ �~$�F0�F4�~L��=�FD_�F<    ��^]� _3�^]� ��������������U��ES�]V���F<    �F@����   ��<tzWS�ND�@������ESPSW�� ���F@��F<u�N�9�V �:�N0��N@��u7��u�ǋV�:�N$���+ЋF4Ӊ�N �9 u�V�:�F �     �N0�9�N@_^[]� ����������U��V�1W�y��u�� 3��Miɔ   �;xw��t�����3�;xs��� �E�x_�0^]� �����U��j�hЈd�    P��SVW�'3�P�E�d�    �e����}�E�������v���"�_������������;�s�����+�;�w�4�NQ���E�    ������E�&�E�M�E�@�e�P�E�������E�jË}�u�]��v �r�G��GSP�E�VRP�� ���r�OQ��  ���M�G�  ��w�_��r��� �M�d�    Y_^[��]� �u�~r�VR�U�  ��j �F   �F    j �F �� �������U����US�]V�uW�}2��E��M��E��E�PQRWVS�����+��g�����������i��   ���_^[��]������������U��E�U;�tS�]VW����x�   ���;�u�_^[]�������U��V�uW�};�tS�]S�������Ɣ   ;�u�[_^]�������U��U��v#�ES�]VW��t�   ����J��x��w�_^[]��U��j�h�d�    P��SVW�'3�P�E�d�    �e��u�}3ۉu�]���$    ;}tU�u�u��E�;�tW���e����Ɣ   �]��u�ǔ   �ыu�};�t��$    ��������Ɣ   ;�u�3�SS�� �ƋM�d�    Y_^[��]���V�qP���5���V�P���� ��^�����V��~r�FP�^�  ��3��F   �F�F^�����������U��VW�y��wP�������V�P��� ���Et	W��  ����_^]� ��������U��yr�AV�uQP��������^]� V�u�AQP���p�����^]� ���������U��j�h(�d�    PQV�'3�P�E�d�    ��u������E3ɉM����u�   �u���t���t���E�x�Pr�@���QRP��������ƋM�d�    Y^��]� ����U��U��V�p�d$ �@��u��M+�P�ARPj ���������^]���������������U��Q�M�U�E� �E�P�EQ�MR�UPQR���������]�����U��Q�M�U�E� �E�P�EQ�MR�UPQR��������]�����U��j�ha�d�    P��SVW�'3�P�E�d�    �e��u�}3ۉu�]���$    ;�vL�u�u��E�;�t�EP������O�Ɣ   �]��u�ԋu�};�t���3����Ɣ   ;�u�3�SS�g� �M�d�    Y_^[��]���������������U��V������~$r�FP���  ��3��F$   �F �ΈF�b� �Et	V��  ����^]� �����̃y$r�AÍA���U��V��� ��~$r�FP�e�  ��3��F$   �F �ΈF�� �Et	V�@�  ����^]� ������U��j�h��d�    PQSV�'3�P�E�d�    ��u�3�S�V� �   �F�^�]��^�F8�^4�^$�FT�^P�^@�Fp�^l�^\�EPV�E��d� ���ƋM�d�    Y^[��]� ������������U��j�h�d�    PQSVW�'3�P�E�d�    ��u�V�E�   �� ���~pr�F\P�V�  ��3ۿ   �~p�^l�^\�~Tr�F@P�4�  ���~T�^P�^@�~8r�F$P��  ���~8�^4�^$�~r�FP���  ���~�^�Έ^�E������d� �M�d�    Y_^[��]���V��~r�FP��  ��3��F   �F�F^�����������U��S�]V�����+F;�w��� ����   W�~����v�� �F;�s9�NQW���������vZ�U�FRSP��������~�~r:�F�8 _��^[]� ��uщ~��r�F_�  ��^[]� �F_�  ��^[]� �F�8 _��^[]� �����U��S�]VW�}��9_s�^� ��E+�;�s���M;�uj��W�������Sj ������_��^[]� ���v��� �M�F;�s�FPW�������M��vj�yr/�I�-��u�~��r�F_�  ��^[]� �F_�  ��^[]� ���~�^r���ËUW�Q�NQP�� ���~�~r��; _��^[]� ����������U��USVW���tF�~�F��r����;�r1��r���ȋ^�;�v��r� �MQ+�RV�������_^[]� �}���v��� �F;�s�VRW��������vY�N�^��r.��,��u�~��r�F_�  ��^[]� �F_�  ��^[]� �ËUWRQP�� ���~�~r��; _��^[]� �����U��Q�UV�uW�}�E� �E�P�ER��QPVW�����΃���+΍�_^��]� ����U��V3���j��F�F   P�F�EP�������^]� ��������U��j�h(�d�    P��D�'3ŉE�SVWP�E�d�    �A � 3҉M�;�t'�A �q0� �6�;�s�A0��A ��Q���K  �AL;��=  9Q<uP�{� ������&  ���!  �E�   �U�U�P�U��Q� �������  Pj�M��Y����}�E؃��5  ���u̅�t!�ȃ�s�M�;�w�ȃ�s�M؋U��;�v�� �}�U�E؍Mԃ��t�ȃ�s�M��;�r��� �}�U�E؋ڃ���   ����t�ȃ�s�M�;�w�ȃ�s�M��;�v�� �}�U�E؍Mԃ��t��s�E��;�r�� �}ċO<��R�E�P�E�P�E�P�E�P�E��PV�GDP�҅���   ��~_����   �}���   j�U�R�M���������7���P�E�jP�2� �uӃ��M��L������   �M؉M̋�������u��%����E�9E���   �U�E؃���   ����t!�ȃ�s�M�;�w�ȃ�s�M؋]��;�v�� �U�E؍Mԃ��t��s�E؋U��;�r�� �E�+�Pj �M��5����OLQ�]� ����������M���������M�d�    Y_^[�M�3���� ��]Íu��b����}�M�Q�M���������+���+}ȋ����~�UċBL�M��T�NPR��� ������uӍM��'���������U��V�u��W�x�I �@��u�+�PV�p���_^]� ����������U��SVW�}���    ��t�E9Fw;Fv�� �E�]���G9^w;^v�t� �]����t;�t�`� �O;�t!�F�E �UR�UR�URQPS�w������F��_^[]� ��������U��j�hX�d�    P��,�'3ŉE�SVWP�E�d�    �y< �M���  �yA ��  ��Pj��҃���m  �   3��E� �M�E؉E��E�   ��s�E��@ �E�    �E؋U����    ����   �؉]̅�t!�ȃ�s�M�;�w�ȃ�s�M؋u��;�v�_� �U�E؍Mԃ��t�ȃ�s�M؋u��;�r�9� �U�E؋}����   ����t$�ȃ�s�M�;�w�ȃ�s�M؋]�ˋ]�;�v��� �U�E؍Mԃ��t��s�E؋U��;�r��� �EЋH<��R�E�P�E��SV��DP�҃� t)��t+���M��7  �>  �]؉]������u��i����E��@A �U�E؃���   ����t!�ȃ�s�M�;�w�ȃ�s�M؋}��;�v�H� �U�E؍Mԃ��t�ȃ�s�M؋}��;�r�"� �U�E؋}�+�tv����   ����t!�ȃ�s�M�;�w�ȃ�s�M؋]��;�v��� �U�E؍Mԃ��t��s�E؋U��;�r�� �EЋHLQWjV�O� ��;�u7�U�E؋MЀyA t4�������Wj�M�����������u������u��h����M�����2��
�M�������M�d�    Y_^[�M�3���� ��]������U��V�uW�};�t���������Ɣ   ;�u�_^]� ���������U��Q�UV�uW�}�E� �E�P�ER��QPVW�������i��   ���_^��]� ����U��Q�U�E� �E�P�ER�U��Q�MPQR��������]� ��U��V�u�~r�FP�*�  ��3��F   �F�F^]� ���U��S�]V�u;�t!W�}j�j V����������;�u��_^[]ËE^[]����������U����'3ŉE����M;�tT�PS�XV�p�]��YW�x�X�Y�X�Y�X�Y�X�Q�U��q�q�y�Q�P�p�q�Q�P_�p^�Q[�M�3��E� ��]� ���U��j�h��d�    PQV�'3�P�E�d�    ��u��� 3��N���j��A�A   P�E��A�EP�����ƋM�d�    Y^��]� �������U��EVP����������^]� ����V������~$r�FP��  ��3��F$   �F �F��^�D� ��������������U��j�h��d�    PQV�'3�P�E�d�    ��u��G� 3��N� �j��A�A   P�E��A�EP�;����ƋM�d�    Y^��]� �������U��Q�V�u3�j���R�F   �VP�ΉU��V�������^��]� �������������U��j�hԊd�    P��   SVW�'3�P�E�d�    3ۉ]��}����   9��   j��  �����u3��E�;�t2�M�E�P�Y���P��`����E��E�   �"���j P�λ   �����E�   ���t�����`����]�������t�}�r�M�Q��  ���   �M�d�    Y_^[��]�������V��� ��~$r�FP���  ��3��F$   �F �F��^�t� ��������������U��UV���W�F   �F    �F �x�@��u�+�PR���}���_��^]� �����U��Q�UV�u3��F�F   �E��F�EPRQ���V�����^��]� �������������V��F��t	P� �  ���P�F    �F    �F    � �  ��^������������U��j�h�d�    P��4�'3ŉE�SVWP�E�d�    �]�щUЃ��u3��  �B$���t �B4�0�;�s��B$��Q������  �BL����  �z< uP��P�� �������  ����  �   3��E� �]̉M�E؉E��E�   ��s�E��@ �E�    �E؋U�I ���	  �؉]ȅ�t!�ȃ�s�M�;�w�ȃ�s�M؋u��;�v�?� �U�E؍Mԃ��t�ȃ�s�M؋u��;�r�� �U�E؋}����  ����t$�ȃ�s�M�;�w�ȃ�s�M؋]�ˋ]�;�v��� �U�E؍Mԃ��t��s�E؋U��;�r�� �EЋH<��R�E�P�SV�E�P�E�P�E�P�EЃ�DP�҅���  ���9  �U�E؃��  ����t!�ȃ�s�M�;�w�ȃ�s�M؋}��;�v�@� �U�E؍Mԃ��t�ȃ�s�M؋}��;�r�� �U�E؋}�+�tz����   ����t!�ȃ�s�M�;�w�ȃ�s�M؋]��;�v��� �U�E؍Mԃ��t��s�E؋U��;�r�� �EЋHLQWjV�G� ��;���   �U�E؋M��AA�M�9M�u|�������}� �M�s{j j�s���������]؉]�������u��Q����u�������u��D�����uB�UЋBL�M�PQ���������t�u�M��T������'�Mԃ���E�������M��9����E��M��,�������M�d�    Y_^[�M�3��m� ��]� �����������U���SV��F W�~@98u�}u�~< u�]K��]�~L ��   �g�����tw��u�}t�M�VLQSR�� ����uX�NL�E�PQ�� ����uD�V 9:u�N�9�V �FA�Ή�V0+ȃ�A�
�E�M��U�_�H�ND^�     �P�H[��]� �E���_3�^��H�H�H[��]� �������������U����EV��~L �MW�}�E��M���   ��������t�FL�U�RP�N� ����uk��t�NLjWQ�� ����uT�FL�U�RP�� ����u@�M�V �ND�N@9
u�FAPPQ�������E�M��U��H�ND_�     �P�H^��]�  �E���_��@    �@    �@    ^��]�  �����������U��QSVW�}���    ��t�E9Fw;Fv��� �E�]���G9^w;^v��� �]����t;�t�� �G;�tB�VPRS�����؋F���E���;�t��I ���I����ǔ   ;}�u�E_�^^[��]� ��_^[��]� ����S��V�s3�;�t(W�{;�t�������Ɣ   ;�u�CP���  ��3�_^�C�C�C[����������������SV��3�W��9^Lt�������u3��FLP�C� ����t3��Έ^H�^A�����^L��=��_�^<�ND^[����U��j�hX�d�    PQVW�'3�P�E�d�    ��u��}W�� 3�j��N����GR�A   �QP�U��Q�����ƋM�d�    Y_^��]� �U��j�h8�d�    P��D�'3�P�E�d�    jh ��M��E�   �E�    �E� �����E�P�M��E�    �G���h8��M�Q�E����� ��U��EVP����������^]� ����U��j�hh�d�    P��SVW�'3�P�E�d�    j �M��� �=t> ��=�E�    �]�u+j �M��c� �=t> u�p>@�p>�t>�M��j� �}�5t>�;ps"�H����u�x t��� ;ps�P�4��3�����uN��t���F�E�WP����������uh4��M��`� h���M�Q��� �u��Ή5�=��k��V�\� ���M��E�������� �ƋM�d�    Y_^[��]��������������U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U��j�h��d�    P��   SV�'3�P�E�d�    �E3ۉ]�����   9��   j��  �����u�]���t7�M�E�P����P��\����E��E�   �U����   �F    ���3��M�E�   �1��t�����\����]�������t�}�r�U�R�9�  ���   �M�d�    Y^[��]�U����US�]V�uW�}2��E��M��E��E�PQRWVS�����+�$I�������������    +ȍ�_^[��]��������U��V�uW�};�t*S3ۃ~r�FP��  ���F   �^�^��;�u�[_^]����U��Q�E�V�u3҉j��N��R�A   �QP�U��Q�`�����^��]����������U��j�h�d�    P��SVW�'3�P�E�d�    �e��u�}3ۉu�]���$    ;}tY�u�u��E�;�tj�S�F   �^W�Έ^��������]��u���ǋu�};�t�]V���r�����;�u�3�SS�	� �ƋM�d�    Y_^[��]���������������U��j�h+�d�    P��   �'3�P�E�d�    �E���A�I#���   �} t	j j �� ��t5hp��M��s����E�P�M��E�    ����h���M�Q�E���b� ��t5hX��M��9����U�R�M��E�   �V���h���E�P�E���(� h@���l���������l���Q�M��E�   ����h���U�R�E����� �M�d�    Y��]� �����U��j�hX�d�    PQVW�'3�P�E�d�    ��u��}W�� 3�j��N� ��GR�A   �QP�U��Q�&����ƋM�d�    Y_^��]� �U��EVP����������^]� ����U��QS3�V��WSS�^$�^�^�F  �F   �^�^�^ �.���j��  ����;�t6�� ���� j �M������ �C���s@�C�M���� �~$_^[��]�_�^$^[��]���������������U��j�h��d�    PQV�'3�P�E�d�    ��u��E�    �����P��  ���M�d�    Y^��]�U��j�h��d�    PQVW�'3�P�E�d�    ��u�����~H �E�    t�����~8�E����������t���f��W��  ���N�V� �M�d�    Y_^��]��U��V���u����Et	V�i�  ����^]� ���������������U��j�h��d�    P��SVW�'3�P�E�d�    �E�P�f��P�E�    �����}������E�������t;j �M��M� �G��v	���sH�G�w����֍M�#��R� ��t
��j���Ћ�E�RP���ҋM�d�    Y_^[��]� ���U��V3�W�}��F�F�F;�u_2�^]� ��I�$	v����PW���������    +ύ��F�F_�V�^]� �����������U��j�h��d�    P��   �'3ŉE�SVWP�E�d�    �e��ًC��u3���K+ȸ���������������} �C  �s��+K�������ыM������º"""+Љ�p���;�s�����;��  ����"""+�;�s3���;�s��j W�?����u+s�ȸ������E������P���U������p���+ƍ�RQ���E�    ������p����E�KRPQ�������U��p�������+ƍ��C�MRPQ�������s�K+θ��������������E��t	V���  ����p�������+ύȋM�S����+эЉK�C�  ��p���R��  ��j j ��� ��+M�u��������������¹   ��t����;Esy�}�E��p�������+�����QRP��������K+M��t���P�������C��������+�WP���E�   �����s�[�E��t���R+�SP� ������N�E����+���p�����P���P+�W���W�����p����UQWR�C�������t���P�E�VP��������M�d�    Y_^[�M�3��q� ��]� ���������������U��j�h&�d�    P��<  SVW�'3�P�E�d�    �e���u�F��u3���N+ȸ��g����������ڋ}����  �N+N���g����������¹�Ϻ+�;�s������8;��m  ���躑Ϻ+�;�s3���;�s��j S�ؿ���M+N�E츧�g����������E�i��   E�3Ƀ��M��M��MQWP��������U�E�NRPQ���E�   �.����U�F�M�iҔ   U��E�   RPQ���	����F�N+ȸ��g�������������F�E�������t�NQP���"����VR���  ���E�i۔   i��   ���^�~�F�M�d�    Y_^[��]� �]����u�}�~�M��i��   �PW�������~ �M�i��   �M�iҔ   �R�V����W�z�  ��j j ��� �N+M���g�����������;���   �MQ��L���辻���E�N��i۔   �RQP���E�   ������N+M��L���R���g�����������+��FWP���E��:���^�v�U��L���Q+�VR�E�   �*�������L����   �E�M�i��   �Q�R�U�P����j j ��� �EP����������i��   �^S��+�SP���E�   �E�6����M�USQR�F����������P�E�WP�������������E������M����M�d�    Y_^[��]� ���������U��Q�M�U�E� �E�P�EQ�MR�UPQR���������]�����U��j�hh�d�    P��SVW�'3�P�E�d�    j �M��� �=�= ��=�E�    �]�u+j �M��� �=�= u�p>@�p>��=�M��� �}�5�=�;ps"�H����u�x t�y� ;ps�P�4��3�����uN��t���F�E�WP���������uh4��M���� h���M�Q�`� �u��Ή5�=�Y]��V�ܸ ���M��E������Q� �ƋM�d�    Y_^[��]��������������U��V�uW�};�tS�]j�j S��������;�u�[_^]������U��Q�E�MV�uPQV�E�    ���������^��]����������U��j�ha�d�    P��SVW�'3�P�E�d�    �e��u�}3ۉu�]���$    ;�vZ�u�u��E�;�t�Ej�S�F   �^P�Έ^�����O���]��u�ǋu�};�t�]V��������;�u�3�SS�� �M�d�    Y_^[��]�U��j�h��d�    PQV�'3�P�E�d�    ��j�s�  3Ƀ�;�t�0�3���N�N�N�ƋM�d�    Y^��]��������U��j�h��d�    PQV�'3�P�E�d�    �M��A��P�D
����q����E�    ������F��H�D1�X��M�d�    Y^��]�������������U��EVWP�����������B�����Є�t�G<    _^]� �ωw<跶��_^]� �U���   �'3ŉE�SV�ًCW�   �u�}��{�u��+ȸ��������������;�vH9{v�� �K+K�E�P���������������+�VWP�������_^[�M�3���� ��]�| s]9{v�J� �K���t����M�;Kv�2� �M���M�V��|�����|����������t����M���|���WPQR��t���P���@����M�_^3�[�� ��]�| �������������U��j�h�d�    P��SVW�'3�P�E�d�    ��^�F�}��+ȸ��g������������E�    ;�v79^v�x� �N+N�EP���g�����������+�WSP�������PsN9^v�?� �F��U�E;Fv�*� �E�W�U܉M�R�M�E�������M�P� SQRP�M�Q��������M�E�����赲���M�d�    Y_^[��] �U��E�UP��Q�MQR������]� �U��j�h�d�    PSVW�'3�P�E�d�    ��3�9^L��   �E�M�UPQR谹 ����;���   ���FH�^A�"����O�N0�N4�G�M�F�F�~ �~$�~L��=Q�ΉFD�^<豳��P�]����������B�����Є�t!�M�^<�X���ƋM�d�    Y_^[��]� �Ή~<諳���M�sX���ƋM�d�    Y_^[��]� 3��M�d�    Y_^[��]� �������U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U��j�hY�d�    P��4�'3ŉE�SVWP�E�d�    �e��u�}3ۉủu��E�   �]�]ԉ]��E�;}te�uĉu��E�;�tj�S�E��F   �^P�Έ^����W���E���������ũ�뻋uȋ}�;�t�]V���6�����;�u�3�SS��� �}�r�M�Q�W�  ���ƋM�d�    Y_^[�M�3��&� ��]�������V�qX�������V�P�致 ��^�����V���HW�13��@u�@(��ȋB0�Ѓ��u�   ��I΅�t�Aǃy( u��j P�E���_��^�U��QV��F��t�M�Q�N�VRQP������VR藶  ���P�F    �F    �F    �w�  ��^��]����������������U��VW�y��wX������V�P�谳 ���Et	W�3�  ����_^]� ��������U��j�h��d�    P��SVW�'3�P�E�d�    �e���u��H�D1΅��(  �I,��t������} ��   ��P�L2����   �MQ����8V��P�E�    �;������M���~U����B�L0(�A �8 �E�   t�Q0�: ~� � ���P�҃��u!��H�D1΃��y( u��j P������W���JHu*�E�������H΃y ue��M�d�    Y_^[��]� ��H�L1(����딋M��B��H���x( u�����H�Hu�E������};Ëu��j j �� �A���y( u��j P����2��M�d�    Y_^[��]� ��������U��SVW�}���    ��t�E9Fw;Fv�� �E�]���G9^w;^v�� �]����t;�t�� �O;�t5�F�E �UR�UR�URQPS������V�؋EP�NQRS�3�����(�^��_^[]� ����U��Q�UV�uW�}�E� �E�P�ER��QPVW�i�������    +΍�_^��]� ��U��SV�uW�}��+ϸ�$I�����������    +ȋE�ɋ�+�;�t+ƉE��E��V�0����;�u�_^��[]�����U��j�h��d�    PQV�'3�P�E�d�    ��u��E���Q�D(��t�H�ذ �E�P�E�    ������F�ƋM�d�    Y^��]� ����U���SV��FW�E�9Fv�� �~�;~v��� �M��QSWP�U�R������_^[��]������������U��j�h�d�    P��SVW�'3�P�E�d�    ���}�3��E�9Et����GX`��E��E�   ��Q�X��G��p����5����_j �Ή^(�F,    �����~( �F0u�F����j P���c����F    ��Q���E�   ����»��������CH �CA �ͬ��3��CL��=�C<�KD�ǋM�d�    Y_^[��]� ������U��j�hW�d�    P��SVW�'3�P�E�d�    ���}�3��E�9Et����GP`��E��E�   ��Q�X��G��p����5����_j �Ή^(�F,    �����~( �F0u�F����j P���c����F    ��Q�E�M��PQ���E�   ���������ǋM�d�    Y_^[��]� �U��j�h��d�    P��SVW�'3�P�E�d�    �e���u�   S3�V�M��}�~�����}� �}���   �}��~{��H�L1(�A �8 �]�t�Q0�: ~� � ���P�҃��u	]��@�M;�u.^��H�L1(�Q �: t�A0�8 ~	��I ���B���
+���s�M��E�    �}�M� �~ u����J��΅�tA�y( u��j P�����E���Q�D(�E�������t�H�\� �ƋM�d�    Y_^[��]� ^�M�ˉM��Q�L2(�W����'����M��@��H���x( u�����H�Hu�E�    �/AËu��?���j j �g� ����������������U��j�h��d�    P��SVW�'3�P�E�d�    �e��u3�WV�M܉}��E� �o����}� �}���   ��I�E�P��"O��P�E��(������M���E� �gN���Mj�W�|�����B�0�A�E���~�����r������I(�A �8 t�Q0�: ~� � ���P�҅�v	���uy�M��E�    �}��@ƀ}� �@    u����I΅�t�Aǃy( u��j P�]����E܋�J�D(�E�������t�H被 �ƋM�d�    Y_^[��]ËS���JH�{����MPj�������H�L1(�E�O茺���K����M��B��H���x( u�����H�Hu�E�    ��BËu�&���j j 蜿 �����U��Q�U�E� �E�P�ER�U��Q�MPQR���������]� ��U��Q�M�U�E� �E�P�EQ�MR�UPQR�;�������]�����U��QVW�}��;��W  �G�O+ȸ�$I����������Eu�������_��^��]� �NS�^+˸�$I�����������9MwY�GSP�GP�M����MQ�N�VRQP�����O+O��$I�������������    +ЋF[��_�N��^��]� ��u3���V+ӉU���$I���U��������9Ew+�G��    +э�SQP�M�����F�O�U��PQR�M��t�FPS���.����FP襫  ���O+O��$I�����������P���������t�N�W�GQRP�������F[_��^��]� ������������U��j�h��d�    P��X�'3ŉE�SVWP�E�d�    �e��E��E��F�u���u�E���N+ȸ�$I����������E��}����  �^��+N��$I����������¹I�$	+�;�s������M��;��  ����I�$	+�;�s�E�    �M��ʉM�;�s�E���j Q������]+^�ȸ�$I��������3���ڋU����E��E�R��    �M�+Í�WQ�Ή]��W����U��E�NRPQ���E�   ������E�ߍ�    +Ӎ��V�EQRP���E�   ������^�N+˸�$I��������������t�VRS���H����FP迩  ���E���    +ȋE�����    +ωV���V�F�  �]����u��}�~��    +ƍ�Q�M�W�������~(�U���    +ȍ���    +ƍ�RQ�M������W�:�  ��j j 蕻 +]��$I�����������;���   �M�Q�M��$����E�N��    +��ۍRQP���E�   �����N+M�U�R��$I�����������+��FWP���E������^�v�U�M�Q+�VR�E�   ��������M��   �M��    +��M��Q���R�U�P�����j j ��� �E�P�M��m����F��    +��P���P+�W���E�   �E�������M��UQWR�F�����E�P�E�SP�T������M�艿���M�d�    Y_^[�M�3��ͭ ��]� �����������U��j�h+�d�    PQV�'3�P�E�d�    ��u��E��F�@   �@    �@ ��E�    ��t0PQ������Q���D��t�    �M�d�    Y^��]� �ƋM�d�    Y^��]� ������������U���SV��^W�~��+ϸ�$I�����������u3��3;�v�P� �M���t;�t�>� �M+ϸ�$I������������M�U�EQjRP���j����^;^v�� �6W�M��u��]�������E�M��U�_^��P[��]� �����U���SVW���G��u3���O+ȸ�$I�����������_��+O��$I�����������;�s.�U�E� �M�Q�MR�GPQjS����������__^[��]� 9_v�R� �U�RSP�E�P������_^[��]� ���������������U��j�h`�d�    PW�'3�P�E�d�    �}�E�E�   ;E,tP��u�� �ML�EP�����E��u�ѷ �E��t#�MQP�y�����J���Dt3��E��E;E,u��}(�UL�r�EP�7�  ���}H�E(   �E$    �E r�M4Q��  ���ǋM�d�    Y_��]���������������U��j�h��d�    P��V�'3�P�E�d�    �ML�UL�E� �E�P�ELQRP�� �̍U,�e�RQ�E�   �������čM�e�QP�E������u��V�E�������T�}(r�UR�e�  ���}H�E(   �E$    �E r�E4P�A�  ���ƋM�d�    Y^��]�������������U�조=��t]��]���������������̡�=���   ��=ǀ�    L�p   �������������������������������U��E�� t��t3�]ù�=��J �����]ø   ]����j j j jdjdhZ� j���G  � ����U��j�h�d�    PQV�'3�P�E�d�    hȪjh�=jH���  ���E��E�    ��t	���   �3�Pj�E������? ��P��=�H�Q`����e�V�ҡ�=�H�Qdj j�h��V�҃�j j�E�   �j? ��PhZ� �E������P ��$�M�d�    Y^��]�����L �����������U��j�hȐd�    PQV�'3�P�E�d�    ��u��L �N�E�    ����]����ƋM�d�    Y^��]������������U��j�hȐd�    PQV�'3�P�E�d�    ��u��N�E�    �x������E������JL �M�d�    Y^��]�����������U��V�������Et	V蹡  ����^]� ��%��%��%��%�������U��E��=� ]�̡�=���   ���   �� Q��Y�������̡�=V��H���   j�V�҃���^����U�존=�UV��H���   RV�Ѓ���^]� �����������U�존=V��H���   j�V�ҡ�=�H�U���   j VR�Ѓ���^]� �����̡�=�P�BQ��Y�U�존=�UV��H���   j VR�Ѓ���^]� ���������U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�EP�EP�EPQ���   �у�]� ���������U�존=VW���H�Qj��ҋ�����u_^]� �U��=�H���   RVW�Ѓ�_��^]� ����������U�존=�P�EPQ�J�у�]� ����U�존=�P�EPQ�J�у����@]� ��������������̡�=�P�BQ��Yá�=�P�BQ�Ѓ����������������U�존=�P�EPQ�J�у�]� ����U�존=�P�EPQ�Jh�у�]� ����U�존=�P�EPQ�Jt�у�]� ����U�존=�P�EPQ�Jl�у�]� ����U�존=�P�EPQ���   �у�]� �U�존=�P�EPQ�Jp�у�]� ����U�존=�P�EPQ���   �у���u]� ��=���   �QP�҃�]� ����U�존=�P�EPQ�J|�у�]� ����U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�EP�EP�EPQ���   �у�]� ���������U�존=�P�EP�EPQ���   �у�]� �������������U�존=�E�P�EQ�$PQ���   �у�]� ����������U�존=�P�E���   ��P�EPQ�M�Q�ҋ�M��P�@�Q�A������]� ���������������U�존=�P�E���   ��0VWP�EPQ�M�Q�ҋ��E���   ���_^��]� ��U�존=�P�EVWP�EPQ���   �ы�=�}���B�H`W�у���t"��=�B�HpWV�ы�=�B�HV�у���_^]� �������������U�존=�P�EVP�EPQ���   �ыu���ΉE��k  �E��tP���n  �UR�{o  ����^]� �U�존=�P�EVWPQ�J\�ы�=�u�����B���   j�V�х�t ��=�B���   j VW�у�_��^]� ��_��^]� ��������������U�존=�P�EPQ�J\�у�]� ����U�존=�P�E���   ��P�EPQ�M�Q�ҋ�M�@�A�������]� �����U�존=�P�EP�EPQ�J$�у�]� U�존=�P�EP�EPQ�J(�у�]� U�존=�P�EP�EP�EPQ���   �у�]� ���������U�존=�E�P�EQ�$PQ�J �у�]� �������������U����E��=�E�   �E��B���   �U�R�URQ�Ћ�=���   �
�E�P�у���]� ������U�존=�P�EP�EPQ�J<�у�]� U�존=�P�EP�EPQ�J@�у�]� U�존=�P�EP�EPQ�J,�у�]� U�존=�P�EP�EPQ�J0�у�]� U�존=�P�EP�EPQ�J8�у�]� U�존=�P�EP�EPQ�J4�у�]� U�존=�P�EPQ���   �у�]� �U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�EP�EP�EPQ���   �у�]� ���������U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�EPQ���   �у�]� �U�존=�P�EPQ���   �ы�=���   �QXP�҃�]� ���������������U�존=�P�EPQ���   �ыU�M��RQ���H ]� ��U�존=�P�EP�EP�EPQ���   �у�]� ���������U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�Eh#  P�EPQ���   �у�]� ��������U�존=�P�EhF  P�EPQ���   �у�]� ��������U�존=�P�EPQ���   �ы�=���   �URP�A`�Ѓ�]� �����������U�존=�P�EPQ���   �у�]� �U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�EP�EPQ���   �у�]� ������������̡�=�P���   Q��Y��������������U��M��U�������Dz"�A�B������Dz�A�B������Dz3�]ø   ]��U����W�E��������u�   �3����U����Az�   �3�3���;���V������Au���]���E�8��$�"� �]���E����E��������z���]���E�8��$�� ���_��^u�E������UF ��_]� ��������������U���V�u�W�}�������Dz�F�G������D{R�G����]�E�$耷 �]�E�F��]�E�$�]��d� �]���E�E�������D{_�   ^��]�_3�^��]�������������U���VW�M������E�}��t-��=�Q4P�B�Ѓ��M��u����_3�^��]Ë�R(���=�H0�QW�҃��M��tԋ�R Q�MQ���ҍM���������t��=�H0���   �U�RW�Ѓ��M�����_��^��]�������������U��VW�}��������=NIVb��   ��   =TCAbgtF=$'  t*=MicM��   j hIicM�������WP�B����_^]� ��BW����_�   ^]� j hdiem��������WP�B����_^]� =INIb��   �~ uŋ�B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� ��  _3�^]� =cnys����_3�^]� ������V���D���=�H0�Vh0[�҉F���F    ��^�����V��F�D���t��=�Q0P�B�Ѓ��F    ^�����̡�=�P0�A���   P�у����������U�존=�P0�E�I���   PQ�҃�]� �������������̡�=�I�P0���   Q�Ѓ���������̡�=�P0�A���   j j j j j j j j j4P�у�(������̡�=�P0�A���   j j j j j j j j j;P�у�(�������U�존=�P0�E�IPQ���   �у�]� ��������������U����E V��P�M������MQh8kds�M�������=�E     �B0���   �M Q�M�U�R�Uj Q�MR�UQ�MR�VQj2R�Ћu ��(�M�������^��]� ������̡�=�I�P0���   Q�Ѓ����������U��V��F��u^]� ��=�Q0�M ���   j j j j j Q�Mj QjP�ҡ�=�H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uË�=�Q0P�B�Ѓ������̋A��u� ��=�Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5�=�v0Q�MQP���   R�U�R�Ћu�    �F    ��=���   j P�BV�Ћ�=���   �
�E�P�у�$��^��]� �������U�존=�P0�E�I�R PQ�҃�]� �U��A��t)��=�Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5�=�v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5�=�v0Q�MQPR�Vl�҃�^]� ����������U��y u3�]� V�u�W�}�؉��ډ��=�P4�A�JlWVP�ы�ډ����ى_^]� �����U��A��u]� ��=�Q4�M�RlQ�MQP�҃�]� ����U��A��u]� ��=�Q4�M�RtQ�MQP�҃�]� ����U��y u3�]� V�u�W�}�؉��ډ��=�P4�A�JtWVP�ы�ډ����ى_^]� �����U���VW��htniv�M������EPhulav�M������hgnlfhtmrf�M�������MQhinim�M������URhixam�M������EPhpets�M������MQhsirt�M������E �}$=  �u�����tPh2nim�M��_���Wh2xam�M��Q����E�U�RP�M�Q���������=���   �Q8P�ҋ�=���   ��U�R�Ѓ��M��L���_��^��]�  ��U���V��htlfv�M������EQ�$hulav�M��&����EPhtmrf�M�������EQ�$hinim�M������EQ�$hixam�M�������EQ�$hpets�M�������M,Qhsirt�M��x��������E ��������Dzn���]$����Dzd�؋U(Rhdauq�M��G����M�E�PQ�U�R���������=���   P�B8�Ћ�=���   �
���E�P�у��M��A�����^��]�( ��Q�$h2nim�M��5����E$Q�$h2xam�M��!����t���������������U����S�]V�EW�}$Wj ���T$���$haerf�E ���\$�E�\$�E�\$��$P�x�������   ��MWj ���T$�$haerf�E ���\$�E�\$�E�\$�C�$Q���3�����tM��UWj ���T$���$haerf�E ���\$�E�\$�E�\$�C�$R�������t_^�   []�  _^3�[]�  ���������U���V��hCITb�M������EPhCITb�M������MQhsirt�M������URhulav�M������M�E�PQ�U�R��������=���   P�B8�Ћ�=���   �
���E�P�у��M�������^��]� ��������U��E��Vj ��P�M�Q�M�u[  �UPR���9�����=�H�Al�U�R�Ѓ���^��]� ����������U��E��UPj ���T$�$htemf�E���\$�E�\$�E�\$�E�$R����]� �����������U��E��Pj ���T$�U�$hrgdf�E���0����(������]�E�\$�E�����]�E�\$�M���]�E�\$�E�$R�%���]� �U��E��Pj ���T$�U�$htcpf�E����������]�E�\$�E���]�E�\$�}�]�E�\$�E�$R�����]� �������������U��Q��u3�]� �E�E�H� V�5�=�v0Q�MQ�M���\$�E�$QPR�V4�҃�^]� ������U��Q��u3�]� �E�H� V�5�=�v0Q�MQPR�V8�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5�=�v0Q�MQPR�V8�҃�^]� ����������U��Q��u3�]� �E�H� V�5�=�v0Q�MQPR�V<�҃�^]� ����������U��SVW���W��t$�E�H�5�=�^0� �uQVP�C<R�Ѓ���u	_^3�[]� �W��t��E�H� ��=�[0Q�NQPR�S<�҃���t̋W��tŋE�H� �=�=�0Q��VP�G<R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5�=�v0Q�MQ�MQPR�VH�҃�^]� ������U��QV3�W��u3��,�E�H� �5�=�v0Q�MQPR�V8��3Ƀ�9M������U�MVR�E�����_^]� �������������U��AV��u3��"�M�Q�	�5�=�v0R�URQP�F8�Ѓ����M�UQ�MR������^]� ��������U��AV��u3��"�M�Q�	�5�=�v0R�URQP�F<�Ѓ����EQ�M�$Q�M������^]� �����U�����V���U��V�U��]�W��t$�E�H� �=�=�0Q�M�QPR�W<�҃���u
_3�^��]� �V��t�E�H� �=�=�0Q�M�QPR�W<�҃���tˋV��tċE�H� �5�=�v0Q�M�QPR�V<�҃���t��M�E�PQ�M�����_�   ^��]� ���U�����A�U�V�U�W�]��u3��&�M�Q�	�5�=�v0R�UR�U�RQP�FH�Ѓ����E�}���t�M�QP���e����E���t�EQ�$P�������_��^��]� ����U��E$�UVP�E��M Q�Mj R�UPQ�Mj R�F���P�EP���:���^]�  �����U��E,�E(�UVj P���\$���E$�M �$Q�E�M���\$�E�\$�E�\$���$R�w����EQ�$P�������^]�( ���U����EVQ�$��MP�H����]��Mj j ���T$�$htemf�E���\$�E�\$�E�\$�E�$Q���w���^]� ��U���E�EVj ���\$���E�M�\$�E�\$���$P�����Q�M�$Q������^]� �����������U���E�EVj ���\$���E�M�\$�E�\$���$P����Q�M�$Q�������^]� �����������U�����V�U�j �U����]���E$�M�\$�E��E �U��\$�E�$PQ�MR�O����M�UP�EPQR������^��]�  ����U�존=�� V��H�A`�U�R�ЋM�E��Qj �U�RP�M�Q�M�����UPR���]�����=�H�Al�U�R�Ћ�=�Q�Jl�E�P�у���^��]� ������������U���HV��M��Q  P�EP�M�Q�M����j j �U�R���S  P�EP���������=�Q�Jl���E�P�у��M��$R  �M��R  ��^��]� ���U�����EV�]���W�}����tQ�$P��������]���M�U��E��U�P�]�Q�U�R��������N��u
_3�^��]� �U�E�r��=�=�0V�uV���\$�E��$P�G4RQ�Ѓ�_^��]� �������������U��E��S�م�u��=�H���   �҅�u[��]� VW��謏  ��htlfv�M�u�j����E�}���]��M�]�E�$諢 �]�E�]��G�$藢 �]���E�M��}��]�E�$hulav����hmrffhtmrf�M��3����}����M�]�E�$�J� �]�E�]�G�$�6� �]���E�M��}�]�E�$hinim�4����}����M�]�E�$��� �]�E�]�G�$�� �]�E�}�]�E���$hixam�M��������Q�$hpets�M������j hdauq�M��s���Vhspff�M��e����E Phsirt�M��T����U�M�QR�E�P���������=���   P�B8�Ћ�=���   �
���E�P�у��M��N���_��^[��]� ���U��E��V���u��=�H���   �҅�u^��]� ���΍  �E�F��u3��"�M�Q�	�5�=�v0R�U�RQP�F<�Ѓ����E���h��M������]�E�\$�M��]�E�$� �����M��@�A��^��]� ����������U����E ��U�]���Vj �]�P��MQ�MR�E�PQ�M�U�R�����MP�EPQ���+���^��]� ����U�����UV�]���E�P�]��ERP������U�M�Q�MR���<�����^��]� ���U��A��u]� �M�Q�	V�5�=�v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� ��=�Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� ��=�Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U�존=�P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� ��=�Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj=P�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5�=�v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M��$ �MQ�U�R�M���$ ��tm�}��E��tN��=���   P�BH�ЋM��I����tQ�W�7��=�[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M��{$ ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5�=�v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� ��=�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� ��=�Q0�M�RTQ�MQ�MQP�҃�]� U��A��u]� ��=�Q0�M�RXQ�MQ�MQ�MQ�MQ�MQP�҃�]� ���̋A��uË�=�Q0P�Bh�Ѓ�������U��A��u]� ��=�Q0�M�R\Q�MQP�҃�]� ����U��A��u]� ��=�Q0�M�R`��   �QP�҃�]� ��U��A��u]� ��=�Q0�M�R`QP�҃�]� ��������U��A��u]� ��=�Q0�M�RdQ�MQ�MQ�MQP�҃�]� ������������U�존=V�u�VW���H4�R�ЋE�F    �~�H� ��=�R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� ��=�Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I��=�R0P�EPQ���   �у�]� ������̡�=�I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u��=� ��=�R0�I�RPV�uVP�EPQ�҃�^]� �����������U�존=�P0�E�I�RtP�EP�EP�EP�EPQ�҃�]� �U�존=�P0�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U��E�P� V�5�=�v0R�UR�UR�UR�URP�A�NxP�у�^]� ��������U��E� ��=�R0j j j j j j j P�A���   jP�у�(]� �����������U��E� ��=�R0j j j j j jj P�A���   jP�у�(]� �����������U��E� ��=�R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M������E�H� ��=�R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R�����M��������^��]� ����������U��E�P� V�5�=�v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5�=�v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5�=�v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5�=�v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U�존=�P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U�존=�UVj j j j j R��H0�E�Vj P���   jR�Ћ�=�Q0�E�N���   PQ�҃�0^]� ���������������U�존=�P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡�=�P0�A���   j j j j j j j j jP�у�(�������U�존=�P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡�=�P0�A���   j j j j j j j j j(P�у�(�������U�존=�P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U�존=�P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡�=�P0�A���   j j j j j j j j jP�у�(������̡�=�P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}�M���tj j���!�����u��tj j���������=�H0�U��B�IpVWP�у�_^[��]� ���������U�존=�P0�E�I���   P�EP�EPQ�҃�]� �����̡�=�P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V���D���=�H0�Vh0[�҉F3��F�F���t��F   ��^�������V��F�D���t��=�Q0P�B�Ѓ��F    ^������U��E�UVj P�E��MQRPj j ���]�����t�~ t
�   ^]� 3�^]� ��U��E�A�I��u3�]� ��=�B0Q�H�у�]� ����U��S�]V�������=ckhc��   tu=cksatY=TCAb��   Wj hdiem�����������PSW���F   �҃~ ��t��t��u3�������P�[���_^��[]� �~ tK��B����^[]� �~ t6���������t+�F    ^�   []� =atnit�MQS������^[]� ^3�[]� ���������U��V��~ ��   W�}����   �$�؈�E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN��=�M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W��  ���F    _^]� �� �.�<�O�^�m�|�����U��V��~ �"  �EW�}�E����   �$�8����E������A��   �   ���E��������   �   ���E��������   �v���E������A��   �b�E������A��uP��������   �E�E��������u3������A{}�,�E���������E������A�����E������DzU����ء�=�U�H0�F���   j j j j j j j RjP���E�U��(R���\$�E�$W蹓  ���F    _^]� �*�A�X�l�������Ή����U���E�E�Uj���\$�E�\$�E�$PR�w���]� ���U���E�E�Uj���\$�E�\$�E�$PR�G���]� ���U���E�E�Uj���\$�E�\$�E�$PR����]� ��̋�3�� ���H�H�H�������������VW��3����9~u��=�H4�V�R�Ѓ��~�~_^����U�존=�P4�E�I�RxPQ�҃�]� �U��U��t3�A��=�I0R���   P�ҋ�=�Q0�M���   QP�҃�]� ��=�P0�E�I���   PQ�҃�]� ���̡�=�P4�A�JP�у������������̡�=�P4�A�JP�у������������̡�=�P4�A�JP�у������������̡�=�P4�A���   P�у���������̡�=�P4�A���   P�у����������U�존=�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U�존=�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U�존=�P4�E�I�R PQ�҃�]� �U�존=�P4�E�I�R$PQ�҃�]� �U�존=�P0�E�I���   P�EP�EP�EPQ�҃�]� ��U�존=�P4�E�I���   PQ�҃�]� ��������������U�존=�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U�존=�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U�존=�P4�E�I�R(PQ�҃�]� �U�존=�P4�E�I�R,P�EP�EPQ�҃�]� ���������U�존=�P4�E�I�R0P�EPQ�҃�]� ������������̡�=�P4�A�J4P��Y��������������U���S�]VW3���~Pj�ˉE�E�����j j�ˉE������E��=�H0�UR�W�E�P�ApR�Ћ�=�Q4�F�JP�ы�=�J0j �U�R�U�R�U�R�U�RP�F�P�AxR�Ѓ�,�} _^[t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ���������U�존=�P4�E�I�R8PQ�҃�]� �U�존=�P4�E�I�R<PQ�҃�]� �U�존=�P4�E�I���   P�EPQ�҃�]� ���������̡�=�P4�A�J@P�у�������������U�존=�P4�E�I�RDP�EPQ�҃�]� �������������U�존=�P4�E�I�RHP�EPQ�҃�]� �������������U�존=�P4�E�I�RLP�EPQ�҃�]� �������������U�존=�P4�E�I�RPP�EPQ�҃�]� �������������U�존=SV�uW�����   �QV�҃�����   ��=���   �]�QS�҃�S��uA��=���   �Q@�ҋء�=���   �Q@V�ҋ�=�Q4�JPSP�GP�у�_^[]� ��=���   �H�у���uD��=���   �H8S�ы�=�؋��   �H@V�ы�=�J4�WSP�AHR�Ѓ�_^[]� hȫh�  螓  ��_^[]� ��=���   �BV�Ѓ�����   ��=���   �]�BS�Ѓ�S��uC��=���   �B@�Ћ�=���   �؋B8V�Ћ�=�Q4�JLSP�GP�у�_^[]� ��=���   �H�у���uD��=���   �H8S�ы�=�؋��   �H8V�ы�=�J4�WSP�ADR�Ѓ�_^[]� hȫh�  詒  ��_^[]� hȫh�  萒  ��_^[]� ������U�존=�P4�E�I��   P�EP�EP�EPQ�҃�]� ��U�존=�P4�E,P�E(P�E$P�E �IP�E�RXP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U�존=�P4�E�I�R\P�EP�EP�EPQ�҃�]� ����̡�=�P4�A�JdP��Y�������������̡�=�P4�A�JhP�у�������������U�존=�P4�E�I���   P�EP�EP�EPQ�҃�]� ��U�존=�P4�E�I�R`P�EP�EP�EP�EP�EPQ�҃�]� �������������U�존=�P4�E�I�RlP�EPQ�҃�]� �������������U��V�uW��t��؉�}��t��ډ��=�P4�A�JlWVP�у���t��ډ��t��ى_^]� �U��V�uW��t��؉�}��t��ډ��=�P4�A�JtWVP�у���t��ډ��t��ى_^]� �U�존=�P4�E�I�RtP�EPQ�҃�]� �������������U���$V��~ ��   ��=�V�H4�AR�Ѓ} t#��=�Q0���   P�F�HQ�҃�^��]� ��hARDb�M܉E��E�    �i���P�M�Q�N�U�R������=���   ��U�R�Ѓ��M�誹��^��]� ���U�존=�P4�E�I�RpPQ�҃��   ]� ������������U�존=�E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U�존=�P4�E�I���   P�EP�EPQ�҃�]� �����̡�=�P4�A���   P�у���������̸   ����������̸   �����������U�존=V��H4�V�A$h�  R�Ћ�=�Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U�존=�P4�E�I�R|P�EP�EP�EPQ�҃�]� �����U�존=�P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}�M���tj j���A�����u��tj j���-������=�H4�U��B�ItVWP�у�_^[��]� ���������U��QSVW�}���3��{���=INIb�   ��   =SACbwt+=$'  t
=MicM�Q  ��P$W����_�   ^��[��]� 3��E��E��@�MQ�U�R���Ѕ�t��=�E�Q4�M�P�FQ�JP�у�_�   ^��[��]� =ARDb��   j j���F���j j�ϋ��9���j j�ωE��+���j j�ωE�����M���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>���p���P���H���P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� j hIicM���T����WP�B ����_^[��]� U�존=�P4�E�I�RXh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M�誴����=�Q4�JpP�FP�у��M������^��]��������V���D���=�H0�Vh0[�҉F���F    ���F   ��^��������V��F�D���t��=�Q0P�B�Ѓ��F    ^������U��VW�}���迵��=cksat`=ckhct�EPW�������_^]� �Fj j j j j j �F   ��=�Q0���   j j j P�у�(��t'_�F    �   ^]� �~ t��B����_^]� _3�^]� �����������U�존=�H��H  ]��������������U�존=�H0���   ]��������������U�존=�H0�U�E��VWRP���   �U�R�Ћ�=�Q�u���B`V�Ћ�=�Q�BpVW�Ћ�=�Q�Jl�E�P�у�_��^��]������������U�존=�H0���   ]��������������U�존=�H0���   ]��������������U��Ej0P�|  ��]��������������U��Ej0P�2�  ��P�Y|  ��]�����U��E�M��j0PQ�U�R�7�  ��P�.|  ��=�H�Al�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P�S�  ��P��{  ��=�Q�Jl�E�P�у���]��U��Ej$P��{  3Ƀ�������]����U��Ej$P�r�  ��P�{  3Ƀ�������]�����������U��E�M��Vj$PQ�U�R�f�  ��P�]{  ��=3Ƀ��B�Pl����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P�r�  ��P�	{  ��=3Ƀ��B�Pl����M�Q�҃���^��]����U�존=�H�U�E��  RPj �у�]���������������U�존=�H�U�ER�UP��  Rj �Ѓ�]�����������U�존=�P4�E�I�R,P�EP�EPQ�҃�]� ���������U�존=�P4�E�I�R0P�EPQ�҃�]� ������������̡�=�P4�A�J4P��Y��������������U���VW�}j ��j������j j�ωE�������E��=�H0�UR�V�E�P�ApR�Ћ�=�Q0�E�H� �RxQ�M�Q�M�Q�M�Q�M�Q�NPQ�҃�(�} _^t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ���U��ESVW�؅�u�Y�}j hdiuM���-�������t3;3u	_^3�[]� j hIicM������;�uj h1icM���Z����uӉ3_^�   []� ��������U���V�uhfnic���J�����tj
��������uShfnic�E�P��蹳���uP�������M��֮�����������t��������uhfnic���#����MQj
���v���^��]��U�존=�P0�E�IP�EP�EP�EPQ���   �у�]� ��U�존=�P0�E�IV�p� ���   V�uj j j V�uVj Pj>Q�҃�(^]� ����U�존=�P0�E�IV�p� ���   V�uV�uj j j�Vj Pj>Q�҃�(^]� ���̡�=�I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V���D���=�H0�WVh0[�ҋ}���F�Ej hmyal���F    �F   �<��F�0����F��t��t�F    j
hhfed�������F_��^]� ���U��VW�}�������=ytsdt�EPW������_^]� ��=�Q0�F���   P�ы�B������_�   ^]� ����������3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ��������������������̸�������������U��E�M� ,  �   �   ]� ��U��Q��=SV��H4�V�AhWR�Ћ�=�Q4�F�JP�ы�=�N�؋B4�PQ�]��ҋV����=�H4�A$h�  R�Ћ�=�Q4�F�JOWKSj j P�ы�=�B4�N�P$h�  Q�ҋN�A<��=�M��X4��0W�%`��To �VP�Cj j R�Ѓ�_^[��]� ����������U���E�Y<]� ���U���V���P(�M�Q���ҋN��t&��=�R0j j j j j j P���   j jQ�Ѓ�(��=�Q�Jl�E�P�ы�=�B�P`�M�Q�ҋF����t ��=�Q0�RXj �M�Qj jj?j P�҃���=�H�Al�U�WR�Ћ�=�Q�J`�E�P�ы�=�B�Pdj j��M�h��Q�ҋF����u3��8��=�E�    �Q0���   �M�Qj j j j j�M�Qh�  jP�ҋ}���(��=�H�Al�U�R�Ѓ���_u3�^��]Ë�=�Q�J`�E�P�ыF����t ��=�J0j �U�Rj j j8j P�AX�Ѓ���=�Q�Jl�E�P�ыF����t��=�J0�Q`jP�҃��F��t���=�E�    �Q0���   �M�Qj j j j j;j h�  jP�҃�(�}� �I����F��t��=�Q0P�Bh�Ѓ��F��t��=�Q0P�Bh�Ѓ��F��t'��=�Q0j j j j j jj j jP���   �Ѓ�(j�M�Q�V(R���E��  �E�    �����������j�v8�v$�q  ���   ^��]����������U���SV��W�~j����  ��V�^<3ۉ^@�^D�^H�^L��=�H0�A h�   R�Ћ�=�Q�J`�E�P�ы�=�B�PdSj��M�h��Q�҃�SS�E�P�M�Q���E��  �]��ֽ����=�B�Pl�M�Q�҃�SSj���V�  _^�C[��]������������̍A�������������U��VW��~D t6�I hȫh�  �a}  j
��z  ��=�HP�V �AR�Ѓ���uC9FDu͋�=�QP�B\�~@W�Ѓ��~D t+hȫh�  �}  ��=�QP�B`W�Ѓ��_3�^]� �M�U�NH�VD��=�HP�Q`�~@W�҃��~D t%�j
�9z  ��=�HP�V �AR�Ѓ���u�9FDu܋�=�QP�B\SW�Ћ^L�FL    ��=�QP�B`W�Ѓ���[_^]� �������U���VW�}����̧��=MicMt<=fnicutj�M�������uP���i����M��Q���jj������_�   ^��]� j hIicM������=���u*j �N(������F�F   ��t��=�Q0P�B�Ѓ��MQW���~���_^��]� ������U��E��V��t3�^]� j�N��  j��n  �F    �v����t��=�H0�QV�҃��   ^]� ��������������j���6�  j�n  ��3�����������U��E3�h�����h  ���P�Ej BR�Uj PR�����]� �U��S�]$V�EW�}�S�]j ����T$���$�E htemf���\$�E�\$�E�\$�E�$P袸������   �G�M�]S��j ���T$�$�E htemf���\$�E�\$�E�\$�E�$Q���W�����t:�E �US���\$���E�\$�E�\$�G�$R�I�����t_^�   []�  _^3�[]�  U���E �ES�]VW�}$W���\$���E�\$�E�\$��$P�K�����th�E �MW���\$�E�\$�E�\$�C�$Q��������t:�E �UW���\$���E�\$�E�\$�C�$R������t_^�   []�  _^3�[]�  ������U���E �ES�]VW�}$W���\$���E�\$�E�\$��$P������th�E �MW���\$�E�\$�E�\$�C�$Q���ݺ����t:�E �UW���\$���E�\$�E�\$�C�$R诺����t_^�   []�  _^3�[]�  ������U��Q�Q��u3���]� �E�H� V�5�=Q�M�Q�E�    �v0PR�VD�ҋ�����t@�E���t9��=�Q�M�RpQP�ҋE�����t��=�QW��P�Bl��W�CC  ��_��^��]� ������U�존=��V��H�A`�U�R�ЋU���M�QR���D�������u��=�H�Al�U�R�Ѓ�3�^��]� �M�Q�M�  ��=�B�Pl�M�Q�҃���^��]� �������U�존=��V��H�A`�U�R�ЋU���M�QR��������M���E�PQ�M�r�����=�B�Pl�M�Q�҃���^��]� ����U���V��M��  �M�E�PQ��� ����M�U���ERP�>����M��  ��^��]� �������������U��EVj ��MP謣���Mh���h  �j j jj PQ��辳��^]� ���������U�����V�U�j �U����]���E$�M�\$�E��E �U��\$�E�$PQ�MR�/����M�UP�EPQR���k���^��]�  ����U�����V�U�j �U����]���E$�M�\$�E��E �U��\$�E�$PQ�MR�ϣ���M�UP�EPQR�������^��]�  ����U�����V�U�j �U����]���E$�M�\$�E��E �U��\$�E�$PQ�MR�o����M�UP�EPQR���;���^��]�  ����U�존=V�uW�����   �QV�҃�V��u,��=���   �Q@�ҋ�=�Q4�J P�GP�у�_^]� ��=���   �H�у���u.��=���   �H8V�ы�=�J4�WP�A$R�Ѓ�_^]� hȫh(  �
u  ��_^]� �U���4��=�H�Q`SVW�}W�ҋu��3�SS�Ή]財��Sj�ΉE�襡����;��   �} ~d��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�h��P�ы�=�B�HW�ы�=�J�U�RP�A0W�Ћ�=�Q�Jl�E�P�у�(��=�B0�M����   VQ�U�R�Ћ�=�Q�J`���E�P�ы�=�B�Pp�M�QV�ҡ�=�H�Al�U�R�Ћ�=�Q�BW�Ћ�=�Q�R0�M�QPW�ҡ�=�H�Al�U�R�Ћu�E��0j ��
S��蕠��j �KQ�ΉE�腠�������������_^[��]���U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj AQj R�UR���-���^]� ��������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR����^]� ����������U��E�E$3҃8��R�U(R�U���\$�E �$R�E���\$�E�\$�E�\$�@�E�$P蒰��]�$ ��������������U��E�@3҃8�]��E��Rj ���T$�$htemf�E���\$�E�\$�E�\$�E�$P�1���]� �������������U��E�E3҃8��R���\$�E�\$�E�\$�@�E�$P�Z���]� ������U��E�E3҃8��R���\$�E�\$�E�\$�@�E�$P芳��]� ������U��E3҃8��R�UR�UR�UR�UP�EPR蔻��]� U��E�E 3҃8��R�U���\$�E�\$�E�$P�EP�ERP�u���]� �U��E�E 3҃8��R�U���\$�E�\$�E�$P�EP�ERP����]� �U��E�E 3҃8��R�U���\$�E�\$�E�$P�EP�ERP����]� �U��E�E 3҃8��R�U���\$�E�\$�E�$P�EP�ERP����]� �U��E3҃8V�u��V��RP�EP����^]� ����������U��Q��u3�]� �E�E�H� V�5�=�v0Q�MQ�M���\$���E�$QPR�V4�҃�^]� ���U��EVj ��MP謜������u�    �F^]� ��u9Ft�   ^]� ���U��EVj ��MP蜜������u�    �F^]� ��u9Ft�   ^]� ���U����EVQ�$��MP�����]����u�E�    �^^]� ��u�F�E������D{�   ^]� ���������������U���$��VW�U����U��M�]�E�PQ�M�U�R觜����x��@�U�}�E����u�V�~_�    �F^��]� ��u�E�P�NQ��������t�   _^��]� ��U�����V���]��M��E��]�PQ�M�U�R�	������@�U��E���u�    �V�F^��]� ��u�E�P�NQ裣������t�   ^��]� ���������������U���VW�}�M�;}u\�uj htsem��������uGPhrdem���ۚ����u6�E�E��EP�M�Q�M�}��^�����t�U�M�R��  _�   ^��]� _3�^��]� �������U���VW�}�M�;}u\�uj htsem���l�����uGPhrdem���[�����u6�E�E��EP�M�Q�M�}��.�����t�U�M�R�^  _�   ^��]� _3�^��]� �������U���SVW�}��;}ua�uj htsem��������uLPhrdem���ۙ����u;��E��E�]P�M�Q�M�}�������t�EQ���$�
  _^�   [��]� _^3�[��]� �U���(�ESW�}�M�;�t;Et	;E��   �]j htsem���\�������   Phrdem���G�����uv�E��M�U��U��U�R�]؉E�M�E�P�M�Q�M�U�R�E�    �E�    �}��E�    �l�����t+�M؋U܃��ĉ�M��P�H�M��z  �   _[��]� _3�[��]� ���U���SVW�}��;}uk�uj htsem��蜘����uVPhrdem��苘����uE��M�E��]���E�P�]�Q�M�U�R�}��c�����t�E��M�PQ���@  _^�   [��]� _^3�[��]� ������̋A���X<Q�ȋB$��j j h����@a  ���������������U�존=��0VW���H�A`�U�R�Ћ�=�Q�J`�E�P�ыE���U�RP�M�Q�M������=�J�U�RP�Ap�Ћ�=�Q�Jl�E�P�ы�=�B�Pl�M�Q�ҡ�=�H�Q`��V�ҡ�=�H�Ap�U�VR�Ѓ����  ��=�Q�Jl�E�P�у�_^��]� ������������U���SVW�}��;}ul�uj htsem��������uWPhrdem���������uF��=�H�A`�U�R�Ѓ��M�Q�M�U�R�}��E�    �����U��u��=�H�AlR�Ѓ�3�_^[��]� ����R��f������  ��=�H�Al�U�R�Ѓ�_^�   [��]� ��U��V�u���B  ��^]� �����������U���<��=SV��H�A`�U�R�Ћ�=�Q�Jd3�Sj��E�h��P���F<�����S�U�SR�E��  �]��XW P�E�P�n�  ��P�M�Q������P�U�R��������=�H�Al�U�R�Ћ�=�Q�Jl�E�P�ы�=�B�Pl�M�Q�҃�9^4tV��=�H4�V0�AR�Ѓ�hARDb�MĉE��]��>���P�M�Q�N4�U�R������=���   ��U�R�Ѓ��M�����9^DtV��=�QP�B\W�~@W�ЋFD��;�t�NHQ�Ѓ��FL�^H�^D�hȫh�  �h  ����=�BP�H`W�у�_^[��]� ������������U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�A�E������D{�   ]� ���������U��V�����u�E�M�U�F�N�    �V^]� ��u�EP�NQ蕛������t�   ^]� ���U��V�����u�E�M�    �F�N^]� ��u�UR�FP�K�������t�   ^]� ���������U��V��~ ���u��=�H4�V�R�Ѓ��E�F    �F    t	V�1  ����^]� �������U��V��F�D���t��=�Q0P�B�Ѓ��E�F    t	V�H1  ����^]� ��������������U���V��3ɍF��H�������=�M��M����   �RQ�M�QP�ҡ�=���   ��U�R�Ѓ���^��]��������������U��V�����u �    ��=�H�Ap���UVR�Ѓ��(��u$��=�Q�R P�EP�NQ�҃���t�   ��=�H�Al�UR�Ѓ�^]� ��U�존=�P�EP�EP�EPQ�Jd�у�]� �����������̡�=V��H$�QDV�҃���^���������U�존=V��H$�QDV�ҡ�=�U�H$�AdRV�Ѓ���^]� U�존=V��H$�QDV�ҡ�=�U�H$�ARV�Ѓ���^]� U�존=V��H$�QDV�ҡ�=�H$�U�ALVR�Ѓ���^]� ��=�P$�BHQ��Y�U�존=�P$�EPQ�JL�у�]� ���̡�=�P$�BQ�Ѓ����������������U�존=�P$�EP�EP�EPQ�J�у�]� ������������U�존=�P$�EP�EP�EPQ�J�у�]� �����������̡�=�P$�BQ�Ѓ����������������U�존=VW�}��H�Q`W�ҡ�=�H$�QV�ҋ�����t ��=�H�QpWV�ҡ�=�H�QV�҃���_^]� ���������U�존=�P$�EPQ�J�у�]� ���̡�=�P$�B(Q��Yá�=�P$�BhQ��Y�U�존=�P$�EPQ�J,�у�]� ����U�존=�P$�EPQ�J0�у�]� ����U�존=�P$�EPQ�J4�у�]� ����U�존=�P$�EPQ�J8�у�]� ����U�존=�UV��H$�ALVR�Ѓ���^]� ��������������U�존=�H$�QDV�uV�ҡ�=�H$�U�ALVR�Ћ�=�E�Q$�J@PV�у���^]���������������U�존=�UV��H$�A@RV�Ѓ���^]� ��������������U�존=�P$�EPQ�J<�у�]� ����U�존=�P$�EPQ�J<�у����@]� ���������������U��V�u���t��=�Q$P�B�Ѓ��    ^]���������U�존=�P$�EP�EPQ�JP�у�]� U�존=�P$�EPQ�JT�у�]� ���̡�=�H$�QX�����U�존=�H$�A\]�����������������U�존=�P$�EP�EP�EPQ�J`�у�]� �����������̡�=�H(�������U�존=�H(�AV�u�R�Ѓ��    ^]��������������U�존=�P(�EP�EP�EP�EP�EP�EPQ�J�у�]� ��=�P(�BQ�Ѓ����������������U�존=�P(�EPQ�J�у�]� ����U�존=�P(�EP�EP�EPQ�J�у�]� ������������U�존=�P(�EP�EPQ�J�у�]� U�존=�P(�EjP�EPQ�J�у�]� ��������������U�존=�P(�EP�EPQ�J�у�]� ��=�P(�B Q�Ѓ���������������̡�=�P(�B$Q�Ѓ���������������̡�=�P(�B(Q�Ѓ����������������U�존=�P(�EPQ�J,�у�]� ����U�존=�P(�EPQ�JP�у�]� ����U�존=�P(�EPQ�JT�у�]� ����U�존=�P(�EPQ�JX�у�]� ����U�존=�P(�EPQ�J\�у�]� ����U�존=�P(�EPQ�J`�у�]� ����U�존=�P(�EPQ�Jp�у�]� ����U�존=�P(�EPQ�Jd�у�]� ����U�존=�P(�EPQ�Jh�у�]� ����U�존=�P(�EPQ�Jl�у�]� ����U�����=V���E�    �E�    �H(�A`�U�RV�Ѓ�����   �E���uI��=�Q�J`�E�P�ы�=�B�M�@pQ�U�R�Ћ�=�Q�Jl�E�P�у��   ^��]� ��=�J��H  h��hH  P�҃��E���u��=�H(�Q,j�V�҃�3�^��]� ��=�Q(�M��Rj QPV�҃���u�E�P��$  ��3�^��]� �M��U�j IQ�MR�e����E�P�$  ���   ^��]� �������������U�존=��V��H�A`�U�R�Ѓ��M�Q������^��u��=�B�Pl�M�Q�҃�3���]� ��=�H$�E�I�U�RP�ы�=�B�Pl�M�Q�҃��   ��]� �U��Q��=�P(�E�PQ�JP�у���u��]� �E3�8U���   ��]� �����U�존=VW�}��H(�QhWV�҃���t$��=�H(�Qh��WV�҃���t_�   ^]� _3�^]� ����U�존=VW�}��H(�QhWV�҃���t>��=�H(�Ah�WRV�Ѓ���t%��=�Q(�Bh��WV�Ѓ���t_�   ^]� _3�^]� ����������U�존=VW�}��H(�QlWV�҃���t>��=�H(�Al�WRV�Ѓ���t%��=�Q(�Bl��WV�Ѓ���t_�   ^]� _3�^]� ����������U��VW�}W��������t8�GP��������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U�존=�P(�EPQ�J0�у�]� ����U�존=�P(�EPQ�J4�у�]� ����U�존=�P(�EPQ�J8�у�]� ����U�존=�P(�EPQ�J<�у�]� ����U�존=�P(�EPQ�J@�у�]� ����U�존=�P(�EP�EPQ�Jt�у�]� U�존=�P(�EPQ�JD�у�]� ����U�존=�E�P(�BHQ�$Q�Ѓ�]� �U�존=�E�P(�BL���$Q�Ѓ�]� ��������������̡�=�H(�Qx�����U�존=�H(�AV�u�R�Ѓ��    ^]��������������U�존=�P(�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J|�у�,]�( ��=�P(�BQ�Ѓ����������������U�존=�P(�EPQ�J�у�]� ����U�존=�P(�EP�EP�EPQ�J�у�]� ������������U�존=�P(�EP�EPQ�J�у�]� U�존=�P(�EjP�EPQ�J�у�]� ��������������U�존=�P(�EP�EPQ�J�у�]� ��=�P(�B Q�Ѓ���������������̡�=�P(�B$Q�Ѓ���������������̡�=�P(�B(Q�Ѓ����������������U�존=�P(�EPQ�J,�у�]� ����U�존=�P(�EPQ�JP�у�]� ����U�존=�P(�EPQ�JT�у�]� ����U�존=�P(�EPQ�JX�у�]� ����U�존=�P(�EPQ�J\�у�]� ����U�존=�P(�EPQ�J`�у�]� ����U�존=�P(�EPQ�Jp�у�]� ����U�존=�P(�EPQ�Jd�у�]� ����U�존=�P(�EPQ�Jh�у�]� ����U�존=�P(�EPQ�Jl�у�]� ����U�����=V���E�    �E�    �H(�A`�U�RV�Ѓ�����   �E���uI��=�Q�J`�E�P�ы�=�B�M�@pQ�U�R�Ћ�=�Q�Jl�E�P�у��   ^��]� ��=�J��H  h��h^  P�҃��E���u��=�H(�Q,j�V�҃�3�^��]� ��=�Q(�M��Rj QPV�҃���u�E�P�  ��3�^��]� �M��U�j IQ�MR�U����E�P�  ���   ^��]� �������������U�존=��V��H�A`�U�R�Ѓ��M�Q������^��u��=�B�Pl�M�Q�҃�3���]� ��=�H$�E�I�U�RP�ы�=�B�Pl�M�Q�҃��   ��]� �U��Q��=�P(�E�PQ�JP�у���u��]� �E3�8U���   ��]� �����U�존=VW�}��H(�QhWV�҃���t$��=�H(�Qh��WV�҃���t_�   ^]� _3�^]� ����U�존=VW�}��H(�QhWV�҃���t>��=�H(�Ah�WRV�Ѓ���t%��=�Q(�Bh��WV�Ѓ���t_�   ^]� _3�^]� ����������U�존=VW�}��H(�QlWV�҃���t>��=�H(�Al�WRV�Ѓ���t%��=�Q(�Bl��WV�Ѓ���t_�   ^]� _3�^]� ����������U��VW�}W��������t8�GP��������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U��VW�}W��� �����t8�GP��������t)�O0Q��������t��HW���������t_�   ^]� _3�^]� ������������U�존=�P(�EPQ�J0�у�]� ����U�존=�P(�EPQ�J4�у�]� ����U�존=�P(�EPQ�J8�у�]� ����U�존=�P(�EPQ�J<�у�]� ����U�존=�P(�EPQ�J@�у�]� ����U�존=�P(�EP�EPQ�Jt�у�]� U�존=�P(�EPQ�JD�у�]� ����U�존=�E�P(�BHQ�$Q�Ѓ�]� �U�존=�E�P(�BL���$Q�Ѓ�]� ���������������U�존=�H(���   ]�������������̡�=�H,�Q����̡�=�P,�B8�����U�존=�H,�A V�u�R�Ѓ��    ^]�������������̡�=�P,�B<�����U�존=�P,�R@��VW�E�P�ҋu����=�H$�QDV�ҡ�=�H$�QLVW�ҡ�=�H$�AH�U�R�Ѓ�_��^��]� �������U�존=�P,�E�RH��VWP�E�P�ҋu����=�H�Q`V�ҡ�=�H�QpVW�ҡ�=�H�Al�U�R�Ѓ�_��^��]� ��̡�=�H,�j j �҃��������������U�존=�P,�EP�EPQ�J�у�]� U�존=�H,�AV�u�R�Ѓ��    ^]�������������̡�=�P,�BQ�Ѓ���������������̡�=�P,�BQ�Ѓ���������������̡�=�P,�BQ�Ѓ���������������̡�=�P,�B,����̡�=�P,�BD����̡�=�P,�B0�����U�존=�P,�R4]�����������������U�존=�H,�A$]�����������������U�존=�H,�AL]�����������������U�존=�H,�A(]�����������������U�존=VW�}��H$�QDW�ҡ�=�H,�QV�ҋ�����t ��=�H$�QLWV�ҡ�=�H$�QV�҃���_^]� ���������U�존=�H�I]�����������������U�존=�H�A]�����������������U�존=�H�I]�����������������U�존=�H�A]�����������������U�존=�H�I]�����������������U�존=�H��\  ]��������������U�존=�H�A ]�����������������U�존=�H�A$]�����������������U�존=�H�I,]�����������������U�존=�H���  ]��������������U�존=�H��p  ]��������������U�존=�H��t  ]��������������U�존=�H��x  ]��������������U�존=�H$�QDVW�}W�ҡ�=�H�Q(���ҋ���t ��=�H$�QLWV�ҡ�=�H$�QV�҃���_^]���������������U�존=�H$�QDVW�}W�ҡ�=�H��X  ���ҋ���t ��=�H$�QLWV�ҡ�=�H$�QV�҃���_^]������������U�존=�H��d  ]��������������U�존=�H�U��L  ��VWR�E�P�ы�=�u���B$�HDV�ы�=�B$�HLVW�ы�=�B$�PH�M�Q�҃�_��^��]����������������U��V�ujV��������^]���������̡�=�H���   ��U�존=�H���   V�uV�҃��    ^]�������������U�존=�P�EP�EP�EPQ���   �у�]� ��������̡�=�P���   Q�Ѓ������������̡�=�P���   Q�Ѓ�������������U�존=�P�EPQ�JL�у�]� ����U�존=�P�EPQ�JP�у�]� ����U�존=�P�EPQ�JT�у�]� ����U�존=�P�EPQ�JX�у�]� ����U�존=�P�EPQ�J\�у�]� ����U�존=�P�EPQ�J`�у�]� ����U�존=�P�EPQ���   �у�]� �U�존=�P�EPQ�Jd�у�]� ����U�존=�P�EPQ�Jh�у�]� ����U�존=�P�EPQ�Jl�у�]� ����U�존=�P�EPQ�Jp�у�]� ����U�존=�P�EPQ�Jt�у�]� ����U�존=�P�EPQ�Jx�у�]� ����U�존=�P�EPQ�J|�у�]� ����U�존=�P�EPQ���   �у�]� �U�존=�P�EPQ���   �у�]� �U�존=�P�EPQ���   �у�]� �U�존=�P�EPQ���   �у�]� �U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�EPQ���   �у�]� �U��E��t ��=�R P�B(Q�Ѓ���t	�   ]� 3�]� U�존=�P �E�RhQ�MPQ�҃�]� U��E��u]� ��=�R P�B,Q�Ѓ��   ]� ������U�존=�P�EPQ�
�у�]� �����U�존=�P�EPQ�J�у�]� ����U�존=�P�EPQ�J�у�]� ����U�존=�P�EPQ�J�у�]� ����U�존=�P�EPQ�J�у�]� ����U�존=�P�EPQ�J�у�]� ����U�존=�P�EP�EPQ���   �у�]� �������������U�존=�E�P�BQ�$Q�Ѓ�]� �U�존=�E�P�B���$Q�Ѓ�]� ���������������U�존=�P�EPQ�J �у�]� ����U�존=�P�EPQ�J$�у�]� ����U�존=�P�EPQ�J(�у�]� ����U�존=�P�EPQ�J,�у�]� ����U�존=�P�EPQ�J0�у�]� ����U�존=�P�EPQ�J4�у�]� ����U�존=�P�EPQ�J8�у�]� ����U�존=�P�EPQ�J<�у�]� ����U�존=�P�EP�EP�EP�EPQ���   �у�]� �����U�존=�P�EPQ�JD�у�]� ����U�존=�P�EPQ���   �у�]� �U�존=�P�EP�EPQ�JH�у�]� ��=�P���   Q�Ѓ�������������U�존=�P�EPQ���   �у�]� �U�존=�P�EPQ���   �у�]� �U�존=�P�EPQ���   �у�]� �U�존=�P�EP�EPQ���   �у�]� ������������̡�=�P���   Q�Ѓ�������������U�존=�P�EP�EPQ���   �у�]� ������������̡�=�P���   Q�Ѓ������������̡�=�P���   Q�Ѓ������������̡�=�P���   Q�Ѓ�������������U�존=�H���   ]��������������U�존=�H���   ]��������������U�존=�H�U�E��VWRP��4  �U�R�Ћ�=�Q�u���B`V�Ћ�=�Q�BpVW�Ћ�=�Q�Jl�E�P�у�_��^��]������������U�존=�H��8  ]��������������U�존=VW�}��H$�QDW�ҡ�=�H$�Q V�ҋ�����t ��=�H$�QLWV�ҡ�=�H$�QV�҃���_^]� ���������U�존=VW�}��H$�QDW�ҡ�=�H$�Q$V�ҋ�����t ��=�H$�QLWV�ҡ�=�H$�QV�҃���_^]� ���������U���V�uV�E�P������������=�Q$�JH�E�P�у���^��]� �������U�존=�P(�} ����PQ�J0�у�]� �������������U�존=VW�}���H(�]�E�QHQ�$V�҃���t-�G��=�H(�]�E�QHQ�$V�҃���t_�   ^]� _3�^]� U�존=VW�}���H(�]�E�QHQ�$V�҃���tO�G��=�H(�]�E�QHQ�$V�҃���t-�G��=�H(�]�E�QHQ�$V�҃���t_�   ^]� _3�^]� ��������������U�존=VW�}���H(�QL���$V�҃���tG��=�G�H(�QL���$V�҃���t)��=�G�H(�QL���$V�҃���t_�   ^]� _3�^]� ����������U��VW�}W���������t8�GP���������t)�OQ���������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W��������t8�GP��������t)�O0Q���������t��HW���������t_�   ^]� _3�^]� ������������U�존=S�]VW���H�QPj S�ҋ�=�H��H  h��Fh�  V�҃��E��u��=�H(�Q,j�W�҃�_^3�[]� ��=�Qj VP�BTS�Ћ�=�Q(�B@VW�Ѓ���t"��=�E�Q(�JVPW�у���t�   �3��UR�Z  ��_��^[]� ��������������U���V�E���MP����P��������=�Q�Jl���E�P�у���^��]� ���U�존=�P(�} ����PQ�J0�у�]� �������������U�존=VW�}���H(�]�E�QHQ�$V�҃���t-�G��=�H(�]�E�QHQ�$V�҃���t_�   ^]� _3�^]� U�존=VW�}���H(�]�E�QHQ�$V�҃���tO�G��=�H(�]�E�QHQ�$V�҃���t-�G��=�H(�]�E�QHQ�$V�҃���t_�   ^]� _3�^]� ��������������U�존=VW�}���H(�QL���$V�҃���tG��=�G�H(�QL���$V�҃���t)��=�G�H(�QL���$V�҃���t_�   ^]� _3�^]� ����������U��VW�}W���������t8�GP���������t)�OQ���������t��$W��������t_�   ^]� _3�^]� ������������U��VW�}W��������t8�GP��������t)�O0Q���������t��HW���������t_�   ^]� _3�^]� ������������U�존=S�]VW���H�QPj S�ҋ�=�H��H  h��Fh�  V�҃��E��u��=�H(�Q,j�W�҃�_^3�[]� ��=�Qj VP�BTS�Ћ�=�Q(�B@VW�Ѓ���t"��=�E�Q(�JVPW�у���t�   �3��UR��  ��_��^[]� ��������������U���V�E���MP�+���P��������=�Q�Jl���E�P�у���^��]� ���U���V�u�E�P��������=�Q$�J�E�P�у���u��=�B$�PH�M�Q�҃�3�^��]á�=�H�A�U�jR�Ѓ���u�M�Q��������t���=�H�QjV�҃���u0��=�H�Q V�҃���u��=�H$�AH�U�R�Ѓ�3�^��]Ë�=�Q$�JH�E�P�у��   ^��]�������U���<��=SVW�E�    ��t�E�P�   ���������=�Q$�JD�E�P�   �у��u���=�B$�}�HDW�ы�=�B$�HLWV�у���t��=�B$�PH�M�Q����҃���t��=�H$�AH�U�R�Ѓ���_^[��]����U��V�u���t��=�QP�B�Ѓ��    ^]���������U��E��t��=�QP���  �Ѓ�]����������������U�존=�H��  ]��������������U�존=�H���  ]�������������̡�=�H���  ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�& ������u_^]Ã} tWj V� ��_������F��=   ^]���U���=�E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�& ������u_^]�Wj V�6 ��_������F��=   ^]�������������U���=�E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�% ������u_^]�Wj V�
 ��_������F��=   ^]�������������U���=�E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�% ������u_^]�Wj V�6
 ��_������F��=   ^]�������������U���=�E��t��s�   �I��H  j j P�҃�]Ã�s�   VW�xW�$ ������u_^]�Wj V�	 ��_������F��=   ^]�������������U��M��t.�=�= t�y���A�uP� ��]á�=�P�BQ�Ѓ�]�������U��M��t.�=�= t�y���A�uP�Q ��]á�=�P�BQ�Ѓ�]�������U�존=�H�U�AR�Ѓ�]��������U�존=�H�U�AR�Ѓ�]��������U���=�E��t#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   VW�xW�B# ������u_^]�Wj V�r ��_������F��=   ^]���������U���=�E��tL�} t#��s�   �U�IR�URP��H  �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   ��=��t�U�IR�URP��H  �Ѓ�]Ã�s�   VW�xW�S" ������u_^]�Wj V� ��_������F��=   ^]����������U��E��w�   ��=��t,�} �U�IR�URPt��H  �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW��! ������u_^]�Wj V�� ��_������F��=   ^]�������U�존=�H�U�AR�Ѓ�]��������U�존=�H�U�AR�Ѓ�]��������U�존=�H�U�AR�Ѓ�]��������U�존=�H�U�AR�Ѓ�]��������U�존=�H|�]�ࡴ=�H|�h   �҃�������������U��V�u���t��=�Q|P�B�Ѓ��    ^]���������U�존=�P|�EP�EPQ�J�у�]� U�존=�P|�EP�EPQ�J�у�]� U�존=�P|�EP�EPQ�J�у�]� U�존=�P|�EPQ�J�у�]� ���̡�=�HL��8  ��U�존=�H@�AHV�u�R�Ѓ��    ^]�������������̡�=�HL�������U�존=�H@�AHV�u�R�Ѓ��    ^]�������������̡�=�PL���   Q�Ѓ�������������U�존=�PL�EP�EPQ���   �у�]� �������������U�존=V��HL���   V�҃���u��=�U�HL���   j RV�Ѓ�^]� ��=���   �ȋBP�Ћ�=���   �MP�BH��^]� �����̡�=�PL��p  Q�Ѓ�������������U�존=�PL�EP�EPQ��t  �у�]� ������������̡�=�HL�Q�����U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U��V�uW�����X����=�U�HL�AVRW�Ѓ�_��^]� �U�존=�PL�EPQ��   �у�]� �U�존=�PL�EP�EPQ�J�у�]� ��=�PL�B Q�Ѓ���������������̡�=�PL�B$Q�Ѓ���������������̡�=�PL�B(Q�Ѓ����������������U�존=�PL�EP�EPQ�J,�у�]� U�존=�PL�EPQ��|  �у�]� �U�존=�PL�EP�EP�EPQ�J0�у�]� ������������U�존=�PL�EP�EP�EP�EPQ�J4�у�]� �������̡�=�PL�B8Q�Ѓ���������������̡�=�PL�B<Q�Ѓ����������������U�존=�PL�EP�EPQ��`  �у�]� ������������̡�=�PL���   Q�Ѓ�������������U�존=�PL��VQ��   �E�P�ыu��P����V���M��W����^��]� �����U�존=�PL�E��T  ��VPQ�M�Q�ҋu��P���V���M���V����^��]� ̡�=�PL�B@Q�Ѓ���������������̡�=�PL�BDj Q�Ѓ��������������U�존=�PL���   ]��������������U�존=�PL���   ]��������������U�존=�PL��4  ]��������������U�존=�PL���   ]��������������U�존=�PL���   ]��������������U�존=�PL��  ]��������������U�존=�PL���   ]��������������U�존=�PL���   ]��������������U�존=�PL��0  ]��������������U�존=�PL�EPQ�JT�у�]� ���̡�=�PL�BQ��Y�U�존=�PL�EP�EPQ�JX�у�]� U�존=�PL�Ej PQ�J\�у�]� ��U�존=�PL�Ej PQ�J`�у�]� ��U�존=�PL�EjPQ�J\�у�]� ��U�존=�PL�EjPQ�J`�у�]� ��U���SVW3��E��P�M��}��}��E��  �}�}���D  W�M�Q�U�R���K  ���M����G7  ��t��=���   ��U�R�Ѓ�_^3�[��]Ë�=���   �J8�E�P�ы�=�����   ��M�Q�҃�_��^[��]��������������U���3�V�E�E�E��P�M��E�   �E�   �E��  �D  j�M�Q�U�R���K  �M��6  ��=���   ��U�R�Ѓ�^��]�����������U�����=�UVW3���}��}����   �I(R�E�P�у��U�R�M��E��  �}�}��C  j�E�P�M�Q���J  �M��6  ��=���   ��M�Q�҃�_^��]� ��U�����=�UVW3���}��}����   �I(R�E�P�у��U�R�M��E��  �}�}��C  j�E�P�M�Q���	J  �M��5  ��=���   ��M�Q�҃�_^��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��B  W�M�Q�U�R���I  ���M����'5  ��t+�u��������=���   ��U�R�Ѓ�_��^[��]� ��=���   �JL�E�P�ыu��P���������=���   ��M�Q�҃�_��^[��]� ���U���SVW3��E��P�M��}��}��E��  �}�}���A  W�M�Q�U�R����H  ���M����g4  ��t+�u���������=���   ��U�R�Ѓ�_��^[��]� ��=���   �JL�E�P�ыu��P���5�����=���   ��M�Q�҃�_��^[��]� ���U���SVW3��E��P�M��}��}��E��  �}�}��4A  W�M�Q�U�R���H  ���M����3  _^��[t��=���   ��U�R�������]Ë�=���   �J<�E�P���]���=���   ��M�Q���E�����]���������������U���SVW3��E��P�M��}��}��E��  �}�}��@  W�M�Q�U�R���TG  ���M�����2  ��t��=���   ��U�R�Ѓ�_^3�[��]Ë�=���   �J8�E�P�ы�=�����   ��M�Q�҃�_��^[��]��������������U���SVW3��E��P�M��}��}��E��  �}�}���?  W�M�Q�U�R���F  ���M����G2  ��t-��u��=����   ���^�U�R�Ѓ�_��^[��]� ��=���   �JP�E�P�ы�@�u��=����   �
�F�E�P�у�_��^[��]� �̡�=�PL��  Q��Y��������������U�존=�PL�E��  ��jPQ�M�Q�ҋ�M�@�A�������]� �������U�존=�PL�E��  ��j PQ�M�Q�ҋ�M�@�A�������]� �������U���SVW3��E��P�M��}��}��E��  �}�}��t>  W�M�Q�U�R���DE  ���M�����0  ��t-��u��=����   ���^�U�R�Ѓ�_��^[��]� ��=���   �JP�E�P�ы�@�u��=����   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��=  W�M�Q�U�R���D  ���M����'0  ��t-��u��=����   ���^�U�R�Ѓ�_��^[��]� ��=���   �JP�E�P�ы�@�u��=����   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}���<  W�M�Q�U�R����C  ���M����g/  ��t-��u��=����   ���^�U�R�Ѓ�_��^[��]� ��=���   �JP�E�P�ы�@�u��=����   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��4<  W�M�Q�U�R���C  ���M����.  ��t��=���   ��U�R�Ѓ�_^3�[��]Ë�=���   �J8�E�P�ы�=�����   ��M�Q�҃�_��^[��]��������������U����E3�V�]��E�E�E��P�M��E�   �E��  �;  j�M�Q�U�R���nB  �M���-  ��=���   ��U�R�Ѓ�^��]� ���������U����EV��M�E�3�Q�M��E�   �E��  �E�E��;  j�U�R�E�P����A  �M��-  ��=���   �
�E�P�у�^��]� ��������U�����=�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��:  j�E�P�M�Q���yA  �M��-  ��=���   ��M�Q�҃�_^��]� ��U�����=�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��
:  j�E�P�M�Q����@  �M��,  ��=���   ��M�Q�҃�_^��]� ��U�����=�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��9  j�E�P�M�Q���y@  �M��,  ��=���   ��M�Q�҃�_^��]� ��U�����=�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}��
9  j�E�P�M�Q����?  �M��+  ��=���   ��M�Q�҃�_^��]� ��U����EV��M�E�3�Q�M��E�   �E��  �E�E��8  j�U�R�E�P���?  �M��+  ��=���   �
�E�P�у�^��]� ��������U���SVW3��E��P�M��}��}��E��  �}�}��48  W�M�Q�U�R���?  ���M����*  ��t-��u��=����   ���^�U�R�Ѓ�_��^[��]� ��=���   �JP�E�P�ы�@�u��=����   �
�F�E�P�у�_��^[��]� ��U���SVW3��E��P�M��}��}��E��  �}�}��t7  W�M�Q�U�R���D>  ���M�����)  ��t��=���   ��U�R�Ѓ�_^3�[��]Ë�=���   �J8�E�P�ы�=�����   ��M�Q�҃�_��^[��]��������������U���SVW3��E��P�M��}��}��E��  �}�}���6  W�M�Q�U�R���=  ���M����7)  ��t��=���   ��U�R�Ѓ�_^3�[��]Ë�=���   �J8�E�P�ы�=�����   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U�����=�UVW3���}��}����   �I,R�E�P�у��U�R�M��E��  �}�}���5  j�E�P�M�Q����<  �M��Q(  ��=���   ��M�Q�҃�_^��]� ��U����EV��M�E�3�Q�M��E�   �E��  �E�E��o5  j�U�R�E�P���^<  �M���'  ��=���   �
�E�P�у�^��]� ��������U����EV��M�E�3�Q�M��E�   �E��  �E�E���4  j�U�R�E�P����;  �M��v'  ��=���   �
�E�P�у�^��]� ��������U�존=�H���   ]��������������U�존=�H���   ]�������������̡�=�H���   �⡴=�H���   ��U�존=�H���   V�u�R�Ѓ��    ^]�����������U�존=�H���   ]��������������U�존=�HL�QV�ҋ���u^]á�=�H�U�ER�UP��@  RV�Ѓ���u��=�Q@�BHV�Ѓ�3���^]����������U�존=�H�U�E��@  R�U�� P�ERP�у�]������U�존=�H���   ]��������������U�존=�H�U �Ej j j j R�Uj P�ER�UP�ER�UP���   R�Ѓ�0]��̡�=�PL�BdQ�Ѓ���������������̡�=�PL�BhQ�Ѓ����������������U�존=�PL�EP�EPQ�Jl�у�]� U�존=�PL�EPQ��d  �у�]� �U�존=�PL�EPQ��  �у�]� ̡�=�PL�BtQ�Ѓ����������������U�존=�PL�EP�EP�EPQ���   �у�]� ���������U�존=�PL�EP�EP�EPQ�J|�у�]� ������������U���<��=SV��HL�QW�ҋ�3ۉ}�;��w  �M���@���M�E�Qh]  �ȉ]ȉ]Љ]ԉ]؉]��E�   �]��}ĉE���F����=���   �PSSW���҅���   ��=�HL�Q W�ҋ���;���   ��    ��=���   �B(���ЍM�Qh�   ���u��;  ������   �M�;���   ��=���   ���   S��;�tm��=���   �ȋB<V�Ћ�=���   ���   �E�P�у�;�t��=�B@�HHV�у���;��]����}��M��?���M��:@����_^[��]� �}���=�B@�HHW�ы�=���   ���   �M�Q�҃��M��J?���M���?��_^3�[��]� ������̡�=�PL���   Q�Ѓ������������̡�=�PL���   Q�Ѓ�������������U�존=�PL�EPQ���   �у�]� ̡�=�PL���  Q�Ѓ������������̡�=�PL���   Q�Ѓ�������������U�존=�PL�EPQ���   �у�]� �U�존=�PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U�E�EVh�h�h�hpR�Q�UR�UR�UQ�A�$�5�=�vLRP���   Q�Ѓ�,^]� ������������̡�=�PL���   Q�Ѓ�������������U�존=�PL�EPQ���   �у�]� �U�존=�PL�EPQ���   �у�]� �U�존=�PL�EPQ���   �у�]� �U�존=�PL�EPQ���   �у�]� �U�존=�PL�EPQ���   �у�]� ̡�=�PL��<  Q�Ѓ�������������U�존=�PL�EP�EP�EPQ��h  �у�]� ���������U�존=�PL���  ]��������������U�존=�PL�EP�EP�EP�EP�EPQ��@  �у�]� �U�존=�PL�EP�EP�EPQ��D  �у�]� ���������U�존=�PL�EP�EP�EP�EPQ��H  �у�]� �����U�존=�HL��$  ]��������������U�존=�HL��(  ]��������������U�존=�HL��,  ]�������������̡�=�HL��\  �⡴=�HL���  ��U���(��=V3��u؉u܉u��u�u�u�u��E�   �u􋈜   ���   W�ҋ}�E�;�t`;�t\��=�QLjP���   ���ЋM��U�Rh=���M�}���  ����=���   ���   �U�R�Ѓ��M؉u��:����_^��]Ë�=���   ���   �E�P�у��M؉u��t:��_�   ^��]����������U���(��=V3��u؉u܉u��u�u�u�u��E�   �u􋈜   ���   W�ҋ}�E�;�t`;�t\��=�QLjP���   ���ЋM��U�Rh<���M�}��	  ����=���   ���   �U�R�Ѓ��M؉u���9����_^��]Ë�=���   ���   �E�P�у��M؉u��9��_�   ^��]����������U�존=�P8�EPQ�JL�у�]� ���̡�=�H8�QD�����U�존=�H8�AHV�u�R�Ѓ��    ^]�������������̡�=�H8�������U�존=�H8�AV�u�R�Ѓ��    ^]��������������U�존=�P8�EP�EP�EPQ�J�у�]� ������������U�존=�P8�EP�EPQ�J �у�]� ��=�P8�B$Q�Ѓ����������������U�존=�P8�EPQ�J(�у�]� ����U�존=�P8�EP�EP�EP�EP�EPQ�J,�у�]� ����U�존=�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U�존=�P8�EP�EPQ�J0�у�]� U�존=�P8�EP�EP�EPQ�J4�у�]� ������������U�존=�P8�EP�EP�EPQ�J�у�]� ������������U�존=�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U�존=�P8�EP�EPQ�J8�у�]� U�존=�P8�EP�EP�EPQ�J<�у�]� ������������U�존=�P8�EPQ�J@�у�]� ����U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H�A0]�����������������U�존=�H�I4]�����������������U�존=�H�Q`V�uV�ҡ�=�H�Q<V�҃���^]�����̡�=�H�Q@�����U�존=�H�ID]����������������̡�=�H�QH����̡�=�H�QL�����U�존=�H�AP]�����������������U�존=�H�AT]�����������������U�존=�H���  ]��������������U�존=�H��|  ]��������������U�존=�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡�=�H���   �⡴=�H��   ��U�존=�H�U�ER�UP�ER�UP���   Rh�,  �Ѓ�]����������������U�존=�H�A]�����������������U�존=�H�Ad]�����������������U�존=�H�Ah]�����������������U�존=�H�Al]����������������̡�=�H�Qp����̡�=�H�Qt����̡�=�H�Qx�����U�존=�H�A|]�����������������U�존=�H���   ]��������������U�존=�H���   ]��������������U�존=�H���  ]��������������U�존=�H��X  ]��������������U�존=�H���   ]��������������U�존=�H���  ]��������������U��V�u��������=�H�U���   VR�Ѓ���^]������U�존=�H���   ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]�������������̡�=�H���   ��U�존=�H���  ]��������������U�존=�H��P  ]��������������U�존=�H��T  ]��������������U��V�u���1����=�H���   V�҃���^]���������̡�=�H���  ��U�존=�H��\  ]��������������U�존=�H�U���   ��R�E�P�ы�M��P�@�Q�A������]�������U�존=�H��  ]��������������U��U�E��=�H�E���   R���\$�E�$P�у�]�U�존=�H���   ]��������������U�존=�H��   ]��������������U�존=�H��h  ]��������������U�존=�H��l  ]��������������U�존=�H��  ]��������������U�존=�H���  ]��������������U�존=�H��$  ]��������������U�존=�H��(  ]��������������U�존=�H��,  ]��������������U�존=�H��0  ]��������������U�존=�H��4  ]��������������U�존=�H��8  ]��������������U�존=�H��<  ]��������������U�존=�H��@  ]��������������U�존=�P���E�P�E�P�E�PQ��D  �у����#E���]����������������U�존=�P���E�P�E�P�E�PQ��D  �у����#E���]����������������U�존=�P���E�P�E�P�E�PQ��D  �у����#E���]����������������U�존=�H���  ]��������������U��V�u(V�u$�E�@��=�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@��=�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U�존=�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U�존=�P0�EP�EP�EP�EPQ���   �у�]� ����̡�=�P0���   Q�Ѓ�������������U�존=�P0�EP�EPQ���   �у�]� �������������U�존=�P0�EP�EP�EP�EPQ���   �у�]� ����̡�=�P0���   Q�Ѓ������������̡�=�H0���   ��U�존=�H0���   V�u�R�Ѓ��    ^]�����������U�존=�H���  ]��������������U�존=�H���  ]�������������̡�=�H���  �⡴=�H��  ��U�존=�H��,  ]��������������U�존=�H��8  ]��������������U�존=�H��0  ]��������������U�존=�H��(  ]��������������U�존=�H��H  ]��������������U�존=�H�U�E���  ��VR�UPR�E�P�ыu�    �F    ��=���   �Qj PV�ҡ�=���   ��U�R�Ѓ� ��^��]��������U���Vj hLGOg�M���*��P�E�hicMCP�k������M��0+����=���   �JT�E�P�у���u(�u���z*����=���   ��M�Q�҃���^��]á�=���   �AT�U�R�Ћu��P���*����=���   �
�E�P�у���^��]�������������U�존=�H��`  ]��������������U�존=�H���  ]��������������U�존=�H�U���  ��V�uVR�E�P�у����S����M��{�����^��]�����U�존=�H���  ]��������������U�존=�H�U���  ��VWR�E�P�ы�=�u���B�H`V�ы�=�B�HpVW�ы�=�B�Pl�M�Q�҃�_��^��]����������������U�존=�H�U���  ��VWR�E�P�ы�=�u���B�H`V�ы�=�B�HpVW�ы�=�B�Pl�M�Q�҃�_��^��]����������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H��   ]��������������U�존=�H��  ]��������������U�존=�H��  ]��������������U��E�M�U��VWPQR�����     �@    ��=���   �M�Rj QP�ҡ�=�H���  �U���R�Ћ�=�Q�u���B`V�Ћ�=�Q�BpVW�Ћ�=�Q�Jl�E�P�у�(_��^��]�����������U�존=�H�U�E��  ��VR�UPR�E�P�ыu�    �F    ��=���   �Qj PV�ҡ�=���   ��U�R�Ѓ� ��^��]��������U�존=�H���  ]��������������U���  �'3ŉE��M�EPQ������R��  ��=�H���  ������Rh���ЋM�3̓���  ��]�������������U�존=�H��h  ��V�U�WR�Ћ�=�Q�u���B`V�Ћ�=�Q�BpVW�Ћ�=�Q�Jl�E�P�у�_��^��]����U�존=�H��l  ��V�U�WR�Ћ�=�Q�u���B`V�Ћ�=�Q�BpVW�Ћ�=�Q�Jl�E�P�у�_��^��]����U�존=�H���  ���҅�tbh���M��%���EPh���M��+���MQh���M��+��j �U�R�E�hicMCP������=���   �
�E�P�у��M��%����]�U�존=�H���  ��V�҅�u��=�H�u�Q`V�҃���^��]�Wh!���M���$���EPh!���M��+��j �M�Q�U�hicMCR�w�����=���   P�BH�Ћ�=�Q�u���B`V�Ћ�=�Q�BpVW�Ћ�=���   �
�E�P�у�$�M���$��_��^��]�����������U�존=�H���  ��V�҅�u��=�H�u�Q`V�҃���^��]�Wh����M��,$���EPh����M��K*��j �M�Q�U�hicMCR������=���   P�BH�Ћ�=�Q�u���B`V�Ћ�=�Q�BpVW�Ћ�=���   �
�E�P�у�$�M��"$��_��^��]�����������U�존=�H���  ���҅�u��]�Vh#���M��t#���EPh#���M��)��j �M�Q�U�hicMCR�������=���   P�B8�Ћ�=���   �
���E�P�у��M��#����^��]������U�존=�H���  ���҅�u��]�Vhs���M���"���EPhs���M��)��j �M�Q�U�hicMCR�_�����=���   P�B8�Ћ�=���   �
���E�P�у��M���"����^��]������U�존=�H��,  ]��������������U�존=�H���  ]��������������U�존=�H��0  ]��������������U��V�u���t��=�QP���  �Ѓ��    ^]������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]�������������̡�=�H���  ��U�존=�H���  ]��������������U�존=�H���  ]�������������̡�=�H���  ��U�존=�H�U���  ��VR�E�P�ыu��P���� ���M��!����^��]�����U�존=�H���  ]��������������U�존=�H��   ]��������������U�존=�H��  ]��������������U�존=�H��  ]��������������U�존=�H��  ]��������������U�존=�H��  ]��������������U���h����M����j �E�P�M�hicMCQ�I�����=���   ��M�Q�҃��M�������]�������U�존=�H��   ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U�존=�H���  ]�������������̡�=�H���  �⡴=�H���  ��U�존=�H��L  ]�������������̡�=�H��P  ��U�존=�H��T  ]������������������������������U�존=�H��|  ]��������������U�존=�H�A`�U��� R�Ћ�=�Q�Jdj j��E�h��P�ыUR�E�P�M�Q��\����=�B�Pl�M�Q�ҡ�=�H�A�U�R�Ћ�=�Q�Jl�E�P�у�,��]��h�=PhD �`v  ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h�=jhD �u  ����t
�@��t]��3�]��������Vh�=j\hD ���\u  ����t�@\��tV�Ѓ���^�����Vh�=j`hD ���,u  ����t�@`��tV�Ѓ�^�������U��Vh�=jdhD ����t  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�=jhhD ���t  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh�=jlhD ���|t  ����t�@l��tV�Ѓ�^�������U��Vh�=h�   hD ���Ft  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�=h�   hD ����s  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�=jphD ���s  ����t�@p��t�MQV�Ѓ�^]� ��=^]� ��U��Vh�=jxhD ���is  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�=jxhD ���)s  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�=jxhD ����r  ����t�@|��t�MVQ�Ѓ����@^]� �   ^]� ������������̋���������������h�=jhD �r  ����t	�@��t��3��������������U��V�u�> t+h�=jhD �Sr  ����t�@��tV�Ѓ��    ^]�������U��VW�}���t0h�=jhD �r  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�=jhD ����q  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�=jhD ���q  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�=j hD ���Lq  ����t�@ ��tV�Ѓ�^�3�^���Vh�=j$hD ���q  ����t�@$��tV�Ѓ�^�3�^���U��Vh�=j(hD ����p  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�=j,hD ���p  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�=j(hD ���Yp  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�=j4hD ���p  ����t�@4��tV�Ѓ�^�3�^���U��Vh�=j8hD ����o  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�=j<hD ���o  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh�=jDhD ���Lo  ����t�@D��tV�Ѓ�^�3�^���U��Vh�=jHhD ���o  ����t�M�PHQV�҃�^]� U��Vh�=jLhD ����n  ����u^]� �M�PLQV�҃�^]� �����������U��Vh�=jPhD ���n  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�=jThD ���ln  ����u^Ë@TV�Ѓ�^���������U��Vh�=jXhD ���9n  ����t�M�PXQV�҃�^]� U��Vh�=h�   hD ���n  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�=h�   hD ���m  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�=h�   hD ���fm  ����u^]� �M���   QV�҃�^]� �����U��Vh�=h�   hD ���&m  ����u^]� �M���   QV�҃�^]� �����U��Vh�=h�   hD ����l  ����u^]� �M���   QV�҃�^]� �����U��Vh�=h�   hD ���l  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh�=h�   hD �el  ����u��=�H�u�Q`V�҃���^��]ËM���   WQ�U�R�Ћ�=�Q�u���B`V�Ћ�=�Q�BpVW�Ћ�=�Q�Jl�E�P�у�_��^��]��U��Vh�=h�   hD ����k  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�=h�   hD ���k  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�=h�   hD ���Fk  ����t���   ��t�MQ����^]� 3�^]� �U��Vh�=h�   hD ���k  ����t���   ��t�MQ����^]� 3�^]� �Vh�=h�   hD ����j  ����t���   ��t��^��3�^����������������U��Vh�=h�   hD ���j  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�=h�   hD ���6j  ����t���   ��t�MQ����^]� ��������U��Vh�=h�   hD ����i  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh�=h�   hD ���i  ����t���   ��t��^��3�^����������������VW��3����$    �h�=jphD �_i  ����t�@p��t	VW�Ѓ����=�8 tF��_��^�������U��SW��3�V��    h�=jphD �i  ����t�@p��t	WS�Ѓ����=�8 tkh�=jphD ��h  ����t�@p��tWS�Ѓ������=h�=jphD �h  ����t�@p��t�MWQ�Ѓ����=�;uG�c����E^��t�8��~=h�=jphD �dh  ����t�@p��t	WS�Ѓ����=�8 u_�   []� _3�[]� U��Vh�=j\hD ���h  ����t3�@\��t,V��h�=jxhD ��g  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�=j\hD ���g  ����t3�@\��t,V��h�=jdhD �g  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�=j\hD ���Vg  ����tG�@\��t@V�ЋEh�=jdhD �E��E�    �E�    � g  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�=j\hD ����f  ����t\�@\��tUV��h�=jdhD �f  ����t�@d��t
�MQV�Ѓ�h�=jhhD �f  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�=j\hD ���If  ������   �@\��t~V��h�=jdhD �#f  ����t�@d��t
�MQV�Ѓ�h�=jhhD ��e  ����t�@h��t
�URV�Ѓ�h�=jhhD ��e  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh�=jthD ���e  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�=j`hD �^e  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh�=���_�����^��]� ������U���Vh�=h�   hD ���e  ����tR���   ��tH�MQ�U�R���ЋuP������h�=j`hD ��d  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t��=���   P�B@��]� �E��t��=���   P�BD��]� ��=���   R�PD��]� �����U�존=�P@���   ]��������������U�존=�P@���   ]��������������U�존=�P@���   ]��������������U�존=�P@���   ]��������������U�존=���   ���   ]�����������U�존=���   ���   ]����������̡�=�P@���   �ࡴ=�P@���   ��U�존=�P@���   ]�������������̡�=�P@���   �ࡴ=���   �Bt��U�존=�P@���   ]�������������̡�=�P@���   ��U�존=�P@���   ]��������������U�존=V��H@�Q$V�ҋM����t��#�����=�Q@P�B V�Ѓ�^]� �̡�=�PH���   Q�Ѓ�������������U�존=�P@�EPQ���   �у�]� ̡�=�P@���   Q�Ѓ������������̡�=�P@�B,Q�Ѓ����������������U�존=�P@�EPQ�J(�у�]� ����U�존=�P@�EP�EP�EPQ�JP�у�]� ������������U�존=�P@�EPQ�JT�у�]� ����U�존=�P@�EP�EPQ�JX�у�]� U�존=�P@�EPQ�J\�у�]� ����U�존=���   �R]��������������U�존=���   �R]��������������U�존=���   �R ]��������������U�존=���   ���   ]�����������U�존=�E���   �E���   P�EP�EQ�$P�EP�EP��]� �����������U�존=���   ���   ]����������̡�=���   �B$�ࡴ=�H@�Ql�����U�존=�H@�Apj�URj �Ѓ�]����U�존=�H@�Apj�URh   @�Ѓ�]�U�존=�H@�U�E�IpRPj �у�]�̡�=���   ����U��V�u���t��=���   P�B�Ѓ��    ^]�����̡�=���   �Q ��U��V�u���t��=���   P�B(�Ѓ��    ^]�����̡�=�H@�Ql�����U��V�u���t��=�Q@P�BH�Ѓ��    ^]���������U�존=�H@���   ]��������������U��V�u���t��=�Q@P�BH�Ѓ��    ^]��������̡�=�PH���   Q�Ѓ�������������U�존=�PH�EPQ���  �у�]� �U�존=�H �Id]�����������������U��}qF u?V�u��t6��=���   �BDW�}W���ЋM��=�B@VQ�HhW�у����w��_^]���̡�=�P@���   ��U�존=�P@���   ]��������������U�존=�P@���   ]�������������̡�=�P@���   ��U��Q��=�P�EWP�M�Q�JP�ы�����u_��]� ��=�B��H  SVh ��_j	S�ы�����u	^[_��]� �M��=�B�U��@TQSVR�Ѓ��> ��^[_��]� ������������U�존=�H�Q`VW�}W�ҡ�=�H�U�ADR�Ћ�����t"��=�Q�BpWV�Ћ�=�Q�BV�Ѓ���_^]���������U�존=�H�Q`V�uV�ҡ�=�H�U�E�I|VRP�у���^]��������������U�존=�H�Q`VW�}W���E��=�H�U�E��R�UP�ERPQ�I@�$�ы�����t"��=�B�HpWV�ы�=�B�HV�у���_^]���U����'3ŉE�V�uW�}�E�0�E�x�   �   ��    ��������
s0�7�D�B��y䡴=�D� �H�Q`W�ҡ�=�H�Adj j��U�RW�ЋM�����_3�^��  ��]�������U��� V�uW�}���&  ��   @vp��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�hX�P�у��U�Rj0j jj �ǋֱ�:�  �U�E�m�P��]�EQ�E��$P�x�������   ����   ��   v`��=�H�A`�U�R�Ћ�=�Q�Jdj j��E�hL�P�у��U�Rj0j jj �ǋֱ
��  �U�E�m�P��]�E�y�����|6��   v,j hH��M������mPj0�P�j jj �]�E�?���j hD��M��e���P�E�WP�
������uPV�@����=�Q�Jl�E�P�ы�=�B�Pl�M�Q�҃�_��^��]���������������U�존=�PT�EP�EPQ�J�у�]� U�존=�PT�EPQ�J8�у�]� ����U�존=�PT�EPQ�J@�у�]� ����U�존=�PT�E�Rh��PQ�M�Q�ҋ�M��P�@�Q�A������]� ������U�존=�HT�U�j R�Ѓ�]�������U�존=�H@�AHV�u�R�Ѓ��    ^]�������������̡�=�HT�j hG  �҃�����������U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U�존=�HT�U�j R�Ѓ�]�������U�존=�H@�AHV�u�R�Ѓ��    ^]�������������̡�=�PD�BQ�Ѓ���������������̡�=�PD�BQ�Ѓ���������������̡�=�PD�BPQ�Ѓ���������������̡�=�PD�BQ�Ѓ���������������̡�=�PD�B(Q�Ѓ����������������U�존=�PX��Q�
�E�P�ы�M��P�@�Q�A������]� �����������U�존=�PX��Q�J�E�P�ы�M��P�@�Q�A������]� ����������U�존=�PX��Q�J�E�P�ы�M��P�@�Q�A������]� ����������U�존=�PX��0VWQ�J�E�P�ы��E���   ���_^��]� �������������U�존=�PX��0VWQ�J�E�P�ы��E���   ���_^��]� �������������U�존=�PX�EPQ�J�у�]� ����U�존=�PX�EPQ�J�у�]� ����U�존=�PX�EPQ�J�у�]� ����U�존=�PX�EPQ�J �у�]� ����U�존=�PX�EPQ�J8�у�]� ����U�존=�PX�EPQ�J(�у�]� ����U�존=�PD�EP�EPQ�J,�у�]� U�존=�HD�U�j j R�Ѓ�]�����U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U�존=�HD�U�j j R�Ѓ�]�����U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U�존=�U�HD�E�	Rj P�у�]���U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U�존=�HD�U�j j R�Ѓ�]�����U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U��U��=�HD�Rj h'  �Ѓ�]��U�존=�H@�AHV�u�R�Ѓ��    ^]�������������̡�=�HD�j j h�  �҃���������U�존=�H@�AHV�u�R�Ѓ��    ^]�������������̡�=�HD�j j h:  �҃���������U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U���3��E��E���=���   �R�E�Pj�����#E���]�̡�=�HD�j j h�F �҃���������U�존=�H@�AHV�u�R�Ѓ��    ^]�������������̡�=�HD�j j h�_ �҃���������U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U��E����u��]� �E���=�E�    ���   �R�E�Pj������؋�]� ̡�=�PD�BLQ�Ѓ����������������U��U��t�M��t�E��tPRQ�`�  ��]������������U�존=�E�PH�B Q�$Q�Ѓ�]� �U�존=�PH�EPQ���   �у�]� �U�존=�PH��0VWQ�JP�E�P�ы��E���   ���_^��]� �������������U�존=�PH��0VWQ�JT�E�P�ы��E���   ���_^��]� �������������U�존=�PH�EPQ���  �у�]� �U�존=�PH�EPQ��   �у�]� �U�존=�PH�EP�EPQ��D  �у�]� �������������U�존=�PH�EP�EPQ��H  �у�]� ������������̡�=�PH���  Q�Ѓ�������������U�존=�PH�EPQ���  �у�]� ̡�=�PH�Bdj Q�Ѓ��������������U�존=�PH�EPj Q�Jh�у�]� �̡�=�PH�BdjQ�Ѓ��������������U�존=�PH�EPjQ�Jh�у�]� �̡�=�PH�BdjQ�Ѓ�������������U�존=�PH�EPjQ�Jh�у�]� ��U�존=�PH�EP�EPQ���   �у�]� �������������U�존=�PH�EP�EPQ���   �у�]� ������������̡�=�PH�BtQ�Ѓ����������������U�존=�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP���P���������t�E��=�QH���   PVW�у���_^]� �����U��EVW���MPQ����������t�M��=�BH���   QVW�҃���_^]� ̡�=�PH��  Q�Ѓ������������̡�=�PH��  Q�Ѓ�������������U�존=�PH�EPQ��  �у�]� �U�존=�PH�EPQ��  �у�]� �U�존=�PH�EP�EPQ��P  �у�]� �������������U�존=�PH�EP�EPQ��  �у�]� ������������̡�=�PH���  Q�Ѓ������������̡�=�PH���  Q�Ѓ������������̡�=�PH���  Q�Ѓ������������̡�=�PH��   Q�Ѓ������������̡�=�PH��$  Q�Ѓ�������������U�존=�PH�EP�EPQ��(  �у�]� �������������U�존=�PH�EP�EP�EPQ��,  �у�]� ���������U�존=�PH�EP�EP�EP�EPQ���  �у�]� �����U�존=�PH�EPQ��<  �у�]� ̡�=�PH��t  Q�Ѓ�������������U�존=�PH�EP�EPQ��@  �у�]� �������������U�존=�PH�EPQ��h  �у�]� ̡�=V��H@�QhWV�҃�j h�  ����������=�HH���   h�  V�҃���
��t_3�^Ë�_^��������������̡�=�P@�BhQ�Ѓ�j h�  �������U�존=�E�PH�E��,  ��P�EPQ�$Q�M�Q�ҋ�M��P�@�Q�A������]� ��������U�존=�E�PH�E��0  ��P�EPQ�$Q�M�Q�ҋ�M��P�@�Q�A������]� ��������U�존=�PH�EP�EPQ��4  �у�]� ������������̡�=�PH��8  Q��Y��������������U�존=�E�PH��<  Q�$Q�Ѓ�]� �������������̡�=�PH��@  Q�Ѓ�������������U�존=�PH�EP�EPQ��D  �у�]� �������������U�존=�E�PH�EP�EQ�$PQ��H  �у�]� �����̡�=�PH���  Q�Ѓ������������̡�=�PH��L  Q�Ѓ������������̋��     �������̡�=�PH����  jP�у���������U�존=�UV��HH���  R��3Ƀ������^��]� ��̡�=�PH����  j P�у��������̡�=�PH��h  Q�Ѓ������������̡�=�PH��l  Q�Ѓ������������̡�=�PH��p  Q�Ѓ�������������U�존=�PH��Q��t  �E�P�ы�M��P�@�Q�A������]� ������̡�=�PH��x  Q�Ѓ�������������U�존=�PH�EPQ��|  �у�]� �U�존=�E�PH���  Q�$Q�Ѓ�]� ��������������U�존=�E�PH���  Q�$Q�Ѓ�]� ��������������U�존=�E�PH���  Q�$Q�Ѓ�]� ��������������U�존=�PH�EPQ���  �у�]� �U�존=�E�HH�U�ER�UP�EQ�$R�UP���   R�Ѓ�]��������������U�존=�E�HH�U�ER�UQ���   �$P�ERP�у�]��U���E�M�`�蜲  �M;�|�M;�~��]�����������U�존=�HH�U�ER�UP���   R�Ѓ�]������������̡�=�PH���   Q��Y�������������̡�=�PH���   Q�Ѓ������������̡�=�PH���   Q��Y��������������U�존=�PH�EP�EPQ���   �у�]� �������������U�존=�PH�EP�EP�EP�EP�EPQ���  �у�]� ̡�=�PH���  Q��Y�������������̋�� l��@    ��l���=�Px�A�JP��Y��������U�존=V��Hx�V�AR�ЋE����u
�   ^]� ��=�Qx�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË�=�QxP�B�Ѓ�������U�존=�Px�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U�존=�E�HH�U�ER�UQ�$P���  R�Ѓ�]������U�존=�HH���  ]��������������U�존=�HH���  ]��������������U�존=�E(�HH�U,�E$R�U Q�$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�(]��������������U�존=�HH���  ]��������������U�존=�E�PH�EPQ�$Q���  �у�]� ����������U���SV���q  �؉]����   �} ��   ��=�HH���  j h�  V�҃��E��u
^��[��]� �MW3��}��  ����   �]��I �E�P�M�Q�MW�O  ��ta�u�;u�Y�I ������u�E�������L�;Ht-��=�Bx�S�@����QR�ЋD������t	�M�P�3  F;u�~��}��MG�}���  ;��v����]�_^��[��]� ^3�[��]� ��������������U�����=SV�ًHH���  j h�  S�]��ҋ�����u
^3�[��]� �E��u��=�HH���  �'��u��=�HH���  ���uš�=�HH���  S�ҋȃ��E��t�W�  ��=�HH���   h�  S3��҃����  ���_�u����    ��=�Hx�U�B�IWP�ы�������   ��=�F�J\�UP�A0R�Ѓ���t�K�Q�M��  ��=�F�J\�UP�A0R�Ѓ���t�K�Q�M�  �E��;Pt&�F��=�Q\�J0P�EP�у���t	�MS�  ��=�v�B\�M�P0VQ�҃���t�M�CP�c  ��=�QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U�존=�HH��  ]�������������̡�=�PH��  Q��Y��������������U�존=�HH���  ]��������������U��Q��V�uW�}Q�$V���&����]��E��E������Au������E������{����]Q�E���$V����_^��]���������U��� ��V�u�U�W�U��}�]�E�PV�M�Q��������E��E�����E��Au���U��������z�����U����E�������z���U�����]���������Au@�����U����E�������z0�����]�U��ER�]�V�E����]��E��]��o���_^��]��]�����������Au����������U�존=�HH�U�j R�Ѓ�]�������U�존=�H@�AHV�u�R�Ѓ��    ^]�������������̡�=�HH�j h�  �҃�����������U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U�존=�HH�Vj h  �ҋ�������   �EPh�  �^�������t]��=�QHj P���   V�ЋMQh(  �4�������t3��=�JH���   j PV�ҡ�=���   �B��j j���Ћ�^]á�=�H@�QHV�҃�3�^]�����U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U�존=�HH�Vj h�  �ҋ�����u^]á�=�HH�U�E��(  RPV�у���u��=�B@�HHV�у�3���^]�����U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U�존=�HH�I]�����������������U�존=�H@�AHV�u�R�Ѓ��    ^]��������������U�존=�PH�EPQ���  �у�]� �U�존=�PH�EPQ���  �у�]� ̡�=�PH���  Q�Ѓ�������������U�존=�HH���  ]��������������U�존=�E�HH�U(�E$R�U P�ER�UP�ER�U���\$�E�$P��p  R�Ѓ�$]������������̡�=�PH��  Q�Ѓ�������������U�존=�PH�EP�EPQ��  �у�]� ������������̡�=�PH��8  Q�Ѓ�������������U�존=�PH�EP�EP�EPQ��   �у�]� ��������̡�=�PH��$  Q�Ѓ������������̡�=�PH��(  Q�Ѓ�������������U�존=�PH�EPQ��0  �у�]� �U�존=�PH�EPQ��4  �у�]� ̋������������������������������̡�=�HH��  ��U�존=�HH��  ]��������������U�존=�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��  �у�0]�, ���������U�존=�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��x  �у�0]�, ���������U�존=�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��  �у�0]�, ���������U�존=�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ��|  �у�0]�, ��������̡�=�PH��X  Q�Ѓ�������������U�존=�PH�EPQ���  �у�]� ̡�=�PH���  Q�Ѓ�������������U�존=�HH��\  ]��������������U�존=�HH��d  ]��������������U�존=��W���HH���   j h�  W�҃��} u�   _��]� Vh�  �����������tq��=�HH���   j VW�҃��M��G����EPh�  �M��f����EQ�$h�  �M��������=�Q@�Jdj �E�PV�у��M�����^�   _��]� ^3�_��]� �����������U��S�]�; VW��u7��=�U�HH���   RW�Ѓ���u��=�QH���   jW�Ѓ���t�   �����   ��=�QH���   W�Ѓ��} u(��=�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;��=�U�HH�ER�USP���  VRW�Ћ�=���   �B(�����Ћ���uŃ; u��=�QH���   W�Ѓ���t3���   �W��u1��=�QH���   �Ћ�=�E�QH���   PW�у�_^[]� ��=�BH���   �у��} u0��=�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ��=�QH�j h  �Ћ؃���u_^[]� ��=���   �u�Bx���Ћ�=���   P�B|���Ѕ�t_���$    ���=�E�QH�MP�Ej Q���  VPW�у���t��=���   �ȋBHS�Ћ�=���   �B(���Ћ���u�_^��[]� ��U��EV���u��=�HH���  �'��u��=�HH���  ���u��=�HH���  V�҃���u3�^]� P�EP������^]� ���������U���H��=�HH���   SV�uWh�  V�ҋء�=�HH�Q|3�Wh�  V�]܉}��҃��E�}�}��}�;��	  ��=���   �B���Ћ�==�  �B  �QH�BxWh:  V�Ћ�=�QH�E䋂�   h�  V�Ћ�=�QHW�؋B|h�  V�]Љ}��Ћ�=�QH�E苂8  V�Ћ�=�QH�E̋�$  V�Ѓ�(�E��E�x���~{�M���M��M̅�tMj�W��M  ���t@�@�Eȃ|� ��~����%�������;�u/����V  ;E�~�E؋��V  E���E��;Pu�E���E��E�G;}�|��}� ts�}�j V�����������  ���x�����tS���-����}�;�uH��=�H��H  �h����h�  S�҃��E���8  �M�SP�,���P��������}ܡ�=�H��H  �h����h�  S�҃��E�����  �M��t��tSQP�;�  ���E؅�~-��=�Qh����h�  P��H  �Ѓ��E�����  ��=�E��QH��(  j�PV�у�����  �}��tjV����������j  �������E���E�    ��=�BH�H|j h�  V��3���9uЉE�u���  �}���}؋��M̅��>  �U�j�R�
L  ����*  �Mȍ@�|� ���]�~����%�������9E��P  ���T  �E�3�3�9C�E܉M���   ��$    �����������tk�]��}������������ϋ9�<��}�@�҉��y�]��|��]�@@�z�<��y�]��|��]�@@�z�<��I�}��]�@���M��}�@����@�M�A;K�M��t����Eԅ���  �+U�j��PR�M��U5  �M�v���E�3�+��U��E��E�9E���   �}� �M����E�t-�M�@���M��U؋U�ʋU؋��U؋R�Q�U؋R�Q;]ԋU��@����M؋M���U؋R�Q�U؋R�Q}b��E��M�9�uU�ыL�����������w4�$�,|�M����4�"�U����t��M����t�
�U����t��;]�|��E��E�F;]������E�;E��z  �U�R�Uu���E�P�Lu���M�Q�Cu����_^3�[��]Ë3�;O�M��Å���   �E�v���W��R�����Q�P�I�H�O��I�M����P�Q���P�I�H��@�E���U�Lv�����P�Q�@�A��t&�G�U�@���U�Lv	�����P�Q�@�A�G��U��@���U�v�����P�Q�@�A�G��w��U��@���U�F�v�����P�Q�@�A��w��U�F�@���U�v�����P�Q�@�A�7F��t+�G�U��@���U�v�����P�Q�@�A�wF���O�E�@��;EЉE��}��N����U�R��s���E�P�s�����  ���   �B����=  ��  ��=�QH�B|j h(  V�Ћ�=�QH�����   h(  V�ЋЃ�3��Uԅ�~!�؋ǅ�t�|� t�K��\K�@;�|�]��]܋�=�Q��H  �[h����h-  S�Ѓ��E�����   �M��t��tSQP���  ���]ԋ�=�Q��H  �h����h2  S�Ѓ��E��tP��t��tSWP赛  ���M����+�=�RH��PQ�E���  V�Ѓ���u�M�Q�r���U�R�xr����_^3�[��]á�=�HH�Q|j h�  V�҉E���=�HH�Q|j h(  V��3�3�3ۃ�9UԉE��}ĉ]���   �u䐋ޅ���   ���E�    ~g�u�<�R��   ����d$ �u��>��\>��EЉY�v�q�u��\7�t7�Y�^���Y�v�]��q�u�B@B����;�|��}ă|� tO�EЋu�8�E��I���R�4����A�F�I�N�M��u���B�R�4����A�F�I�N�u�B<މ}�C;]ԉ]������M�3�3�;�~�U��t���   @;�|�U�R�q�����E�P�q����_^�   [��]ÍI pw{w�w�w����U��E� �M+]� ���������������U��V��V�l���=�Hx�AR�Ѓ��Et	V�s������^]� ����������U�존=�H ���   ]��������������U�존=�H@�AHV�u�R�Ѓ��    ^]�������������̡�=�H �������U��V�u���t��=�Q P�B�Ѓ��    ^]���������U�존=�P �EPQ�JP�у�]� ����U�존=�P �EPQ�J�у�]� ����U�존=�P �EPQ�J�у�]� ���̡�=�P �BQ��Y�U��V�uW�����/�����=�H �Q VW�҃�_��^]� �����U�존=�P �EPQ�J$�у�]� ���̡�=�P �BDQ�Ѓ���������������̡�=�P �BLQ�Ѓ����������������V������̭�F    ��^��������U��E�A�   ]� ��������������U��E�M� P   �P   �   ]� ��� �������������V��W�~���B��3��G�̭��F�F_��^�����������V����t��=�Q P�B4�Ѓ��N^���������������U��E��S�]V��F�K�N��u^[��]�, W�}(�v��tj�U�R�FP�ˉ}��E�    �����K�]0�FS�],��=�R SW�}$W�} W�}W�}W�}W�}WP�FQ�J0P�у�03҅���_�^[��]�, ���U���V��> t6�M��*���hNIVb�M�������=�H ��I8j �U�RP�у��M�����^��]��������U����t*�y t$�y t��=�Q �M�R8Q�MQP�҃�]� 3�]� �������U��V��FW�}��t&���t �x t�x t��=�P �B8jWQ�Ѓ��MQW�����_^]� �������U��V���
���Et	V�o������^]� ��������������̡�=�H\�������U�존=�H\�AV�u�R�Ѓ��    ^]�������������̡�=�P\�BQ��Yá�=�P\�BQ�Ѓ���������������̡�=�P\�BQ�Ѓ����������������U�존=�P\�EPQ�J�у�]� ����U�존=�P\�EP�EPQ�J�у�]� U�존=�P\�EPQ�J�у�]� ���̡�=�P\�B Q�Ѓ����������������U�존=�P\�EPQ�J$�у�]� ����U�존=�P\�EP�EPQ�J(�у�]� U�존=�P\�EP�EP�EPQ�J,�у�]� ������������U�존=�P\�EPQ�J4�у�]� ����U�존=�P\�EPQ�JD�у�]� ����U�존=�P\�EPQ�JH�у�]� ���̡�=�P\�B8Q�Ѓ����������������U�존=�P\�EP�EPQ�J<�у�]� U�존=�P\�EPQ�J@�у�]� ����U���SVW�}��j �ωu��&\����=�H\�QV�҃���S���\��3���~=��I ��=�H\�U�R�U��EP�A,VR�ЋM��Q����[���U�R����[��F;�|�_^[��]� ���������������U���VW�}�E��P���XX���}� ��   ��=�Q\�B V�Ѓ��M�Q���1X���E���t]S3ۅ�~H�I �UR���X���E�P���
X���E;E�!����=�Q\P�BV�ЋE@��;E��E~�C;]�|�[_�   ^��]� _�   ^��]� h�=Ph�f �p#  ���������������U���Vh�=h�   h�f ���C#  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh�=h�   h�f ���"  ����t���   ��t�M�UQ�MRQ����^]� U���Vh�=h�   h�f ���s"  3Ƀ�;�t@���   ;�t6�M�Q���ЋM���P�Q�P�Q�P�Q�P�@�Q�A��^��]� �E�   � �  �P�P�H�H�H^��]� ������U��Vh�=h�   h�f ����!  ����t���   ��t�M�UQ�MRQ����^]� U��Qh�=h�   h�f �!  ����t���   �E���t�EP�U�����]������]�������������U���h�=h�   h�f �V!  3Ƀ�;�tK9��   tC�E���   ���M��$Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]ËE�   � �  �P�P�H�H�H��]��U��h�=h�   h�f ��   ����t���   ��t]��]����U��h�=h�   h�f �   ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h�=h�   h�f �9   ����t���   ��t]���E��M��P�Q�P�Q�P�Q�P�Q�@�A3�]����������U��h�=h�   h�f ��  ����t���   ��t]�����]�U���Vh�=h�   h�f �  ����tZ���   ��tP�M�UWQR�M�Q�Ћ�=�u���B�H`V�ы�=�B�HpVW�ы�=�B�Pl�M�Q�҃�_��^��]á�=�H�u�Q`V�҃���^��]����������h�=h�   h�f �  ����t���   ��t��3��������U��h�=h�   h�f ��  ����t���   ��t]��]����U��M��U+u&�A+Bu�A+Bu�A+Bu�A+Bu�A+B]����������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���E+t��3�����]� �Q+Pu�Q+Pu�Q+PuۋQ+PuӋI+H3�����]� ������U���h�=�   h�   h�f �E��  �E��E��E�    �E�    �E�    �_  ����t���   ��t	�M�Q�Ѓ��UR�E�P��������]��U��E��u��=�MP�EPQ�s�����]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h �j;h�=j�e������t
W���4���3��F��u_^]� �~ t3�9_��^]� ��=�H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ��=�H<�Q��3Ʌ����^��������������̃y t�   ËA��uË�=�R<P��JP�у��������U����u��=�H�]� ��=�J<�URP�A�Ѓ�]� ���������������U���=��u��=�H�]Ë�=�J<�URP�A�Ѓ�]�U���=��$V��u��=�H�1���=�J<�URP�A�Ѓ�����=�Q�J`�E�SP�ы�=�B�Pp�M�QV�ҡ�=�H�A`�U�R�Ћ�=�Q�Jdj j��E�hH�P�ы�=�Bj �M�Q�U�R�P$�M�Q�҅���=�H�Al�U�R���Ѓ�4��[t.��=�Q�u�B`V�Ћ�=�Q�Jl�E�P�у���^��]Ë�=�B�M��@,jQ�U�R�Ћ�=�Q�E�M�PQ�J0�E�P�ы�=�B�u�H`V�ы�=�B�Pp�M�VQ�ҡ�=�H�Al�U�R�Ѓ�(��^��]�U���=��$SV��u��=�H�1���=�J<�URP�A�Ѓ�����=�Q�J`�E�P�ы�=�B�Pp�M�QV�ҡ�=�H�A`�U�R�Ћ�=�Q�Jdj j��E�hH�P�ы�=�Bj �M�Q�U�R�P$�M�Q�҅���=�H�Al�U�R���Ѓ�4��t/��=�Q�u�B`V�Ћ�=�Q�Jl�E�P�у���^[��]Ë�=�B�M��@,jQ�U�R�Ћ�=�Q�E�M�PQ�J0�E�P�ы�=�B�P`�M�Q�ҡ�=�H�Adj j��U�hH�R�Ћ�=�Qj �E�P�M�Q�J$�E�P�ы�=���B�Pl�M�Q���҃�@��t-��=�H�u�Q`V�ҡ�=�H�Al�U�R�Ѓ���^[��]Ë�=�Q�E��R,jP�M�Q�ҡ�=�H�U�E�RP�A0�U�R�Ћ�=�Q�u�B`V�Ћ�=�Q�Jp�E�VP�ы�=�B�Pl�M�Q�҃�(��^[��]�����������U���=��$SV��u��=�H�1���=�J<�URP�A�Ѓ�����=�Q�J`�E�P�ы�=�B�Pp�M�QV�ҡ�=�H�A`�U�R�Ћ�=�Q�Jdj j��E�hH�P�ы�=�Bj �M�Q�U�R�P$�M�Q�҅���=�H�Al�U�R���Ѓ�4��t/��=�Q�u�B`V�Ћ�=�Q�Jl�E�P�у���^[��]Ë�=�B�M��@,jQ�U�R�Ћ�=�Q�E�M�PQ�J0�E�P�ы�=�B�P`�M�Q�ҡ�=�H�Adj j��U�hH�R�Ћ�=�Qj �E�P�M�Q�J$�E�P�ы�=���B�Pl�M�Q���҃�@��t-��=�H�u�Q`V�ҡ�=�H�Al�U�R�Ѓ���^[��]Ë�=�Q�E��R,jP�M�Q�ҡ�=�H�U�E�RP�A0�U�R�Ћ�=�Q�J`�E�P�ы�=�B�Pdj j��M�hH�Q�ҡ�=�Hj �U�R�E�P�A$�U�R�Ћ�=�Q�Jl���E�P���у�@��t/��=�B�u�H`V�ы�=�B�Pl�M�Q�҃���^[��]á�=�H�U��I,jR�E�P�ы�=�B�M�U�QR�P0�M�Q�ҋu���E�P���5�����=�Q�Jl�E�P�у���^[��]���������U���=��$SV��u��=�H�1���=�J<�URP�A�Ѓ�����=�Q�J`�E�P�ы�=�B�Pp�M�QV�ҡ�=�H�A`�U�R�Ћ�=�Q�Jdj j��E�hH�P�ы�=�Bj �M�Q�U�R�P$�M�Q�҅���=�H�Al�U�R���Ѓ�4��t/��=�Q�u�B`V�Ћ�=�Q�Jl�E�P�у���^[��]Ë�=�B�M��@,jQ�U�R�Ћ�=�Q�E�M�PQ�J0�E�P�ы�=�B�P`�M�Q�ҡ�=�H�Adj j��U�hH�R�Ћ�=�Qj �E�P�M�Q�J$�E�P�ы�=���B�Pl�M�Q���҃�@��t-��=�H�u�Q`V�ҡ�=�H�Al�U�R�Ѓ���^[��]Ë�=�Q�E��R,jP�M�Q�ҡ�=�H�U�E�RP�A0�U�R�Ћ�=�Q�J`�E�P�ы�=�B�Pdj j��M�hH�Q�ҡ�=�Hj �U�R�E�P�A$�U�R�Ћ�=�Q�Jl���E�P���у�@��t/��=�B�u�H`V�ы�=�B�Pl�M�Q�҃���^[��]á�=�H�U��I,jR�E�P�ы�=�B�M�U�QR�P0�M�Q�҃�j hH��M���y����=�Hj �U�R�E�P�A$�U�R�Ћ�=�Q�Jl���E�P���у����Q�����=�H�U��I,jR�E�P�ы�=�B�M�U�QR�P0�M�Q�ҋu���E�P���Ջ����=�Q�Jl�E�P�у���^[��]���������U�존=�H<�A]����������������̡�=�H<�Q�����V��~ u>���t��=�Q<P�B�Ѓ��    W�~��t���z)��W��X�����F    _^��������U���V�E�P����T����P���C����M���9)����^��]��̃=�= uK��=��t��=�Q<P�B�Ѓ���=    ��=��tV����(��V�jX������=    ^������������U���8��=�H�A`S�U�V3�R�]��Ћ�=�Q�JdSj��E�hL�P�ы�=�B<�P�M�Q�ҋ�=�H�Al�U�R�Ѓ�;�u^3�[��]�V�M�]���  �M�Q�U�R�M��(  ����   W�}�}���   ��=���   �U��ATR�Ћ�����tF��=�Q�J`�E�P���у��U�Rj�E�P��謺����=�Qj WP�B �Ѓ��E���t�E� ��t��=�Q�Jl�E�P����у���t��=�B�Pl�M�Q����҃��}� u"�E�P�M�Q�M��[  ���7����E�_^[��]ËU��U�_�E�^[��]����������U��E����u��]�VP�M��  �EP�M�Q�M��E�    �E    ��  ����   �u�E���tB��t=��u[��=���   �M�PHQ�ҋ�=�Qj VP�B �Ѓ���u-�   ^��]Ë�=���   �E�JTP��VP�V�������uӍUR�E�P�M��o  ���{���3�^��]�V��~ u>���t��=�Q<P�B�Ѓ��    W�~��t���J&��W��U�����F    _^�������̋�� \����������\����������̅�t��j�����̡�=�P��l  �ࡴ=�P��x  ��U�존=�P��p  ��V�E�P�ҋuP���%���M��%����^��]� ��������̡�=�P��t  ��U�존=�H��d  ]��������������U�존=�H��  ]�������������̡�=�H��h  ��U�존=�H��<  ]��������������U�존=�H���  ]��������������U�존=�H���  ]��������������U���EV���\�t	V�HT������^]� �������������̸   � �������̸   @� �������̸   � �������̸   � ��������U�존=�H�Q`V�uV�҃���^]� �3�� �����������3�� �����������U����   h�   ��@���j P�$]  �M�Eh�   ��@���R�M��MPQjǅ`���    �Y}���� ��]���U����   V�u��u3�^��]�h�   ��@���j P��\  �M�U�Eh�   �M���@���Q�U��U��@����ERPj��`���ǅD������E�`��E����E�p��E����E����E�P��E����|���� ^��]�������������U���   SV�u(3ۉ]���u��=�H�Al�UR�Ѓ�^3�[��]Ë�=�Q�JW�EP3��у����'  �1  �E���tq�UR�M��e"��Wh`��M���q��P�M��N"���u�Wj��E�P�M�Q��\���R�_?�AN����P��x���P�$����P�M�Q�$����P����2  �E���t�E� �� t�M�����L"����t��x�������9"����t��\�������&"����t�M̃���"����t��=�B�Pl�M�Q����҃���t�M���!���}� t"�E(�M$�U�P�EQ�MR�UPQR����������E�P�0  ����M$�U�EVQ�Mj RPQ����������=�B�Pl�MQ�҃���_^[��]�����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`�����������U�존=���   �BXQ�Ѓ���u]� ��=���   �M�RQ�MQP�҃�]� U�존=���   �BXQ�Ѓ���u]� ��=���   �M�R8Q�MQP�҃�]� U��EV��j ���=�Qj j P���   �ЉF����^]� ��=Vj ��H����   j j R�Ѓ��F^�������������U��V��F��u^]� ��=�Q�MP�EP�Q���   P�у��F�   ^]� �U�����W��������Au���]��W���G��Au���]��E��`�������A�  �E����������  ���p�������AuI������AuBV�;r  ���4r  �ȋ��ƙ����ʅ�u�u��E�^�]���E����������__��]�������������Au������=h���������Au>�����]������]������O�_�E��E�����������Au�����U��_�E�������������I �E��E�����x  �]��E��]��E��U��d�����t���E����������__��]���������__��]���������__��]����������������U��M��P]����U��M��P]����U��M��P]����V���|��F    ��=�HP�Q|h��Vh��hp��҉F����^���������̃y �|�u��=�PP�A�JP��Y��U��A��u]� ��=�QP�M�RxQ�MQ�MQP�҃�]� U��A��t��=�QP�M���   QP�҃�]� ���������U��A��t��=�QP�M�RTQP�҃�]� �����������̡�=�HP�Q@�����U�존=�HP�ADV�u�R�Ѓ��    ^]�������������̋��     �@    �V����t)��=�QPP�B<�Ћ�=�QP��J,P�у��    ^�������������U��SV�ً3�W;�t��=�QPP�B,�Ѓ��3�s�}�Eh��W�C��=�QP���   h��hp�P�EP�у�9u�~J���z u!���@   ��=�QP���H�RQ�҃���=�HP��A0VR�Ћ�F��;u�A|�3�9_^��[]� ��������U��SVW��3�9w~<�]��=�HP��A0VR�Ѓ���t-��=�QPj SjP�Bx�Ѓ���tF;w|�_^�   []� ��=�QP��J<P�у�_^3�[]� �����������̡�=�PP��J4P�у�������������̡�=�PP��J8P��Y��������������̡�=�PP��J<P��Y���������������U��U�E�@R�URP�I���]� �����U��V��~ �|�u��=�HP�V�AR�Ѓ��Et	V�.J������^]� ����U��E��u�E�M��=��=�   ]� �����������U��EHV����   �$�X��   ^]á�=@��=��uT�EP�'�����=�,  }�����^]Ëu��t�h��jgh�=j�KJ������t ���M����=��tV�������   ^]���=    �   ^]ËM�UQR腥���������H^]�^]�0����-�=u.�R����m�����=��t�����V�I������=    �   ^]Ã��^]ÍI p�	��h�O��U��E�M�UP��P�EjP�Cw����]��������������̸   �����������U��V�u��t���u6�EjP�Dw������u3�^]Ë��qx����t���t��U3�;P��I#�^]�������U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��5�E��}���t�u+��\�P@�m���u�EH�E����   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}�u�C�]�M��E��VP�҅��c����F��}��t�M�+�I�I �\�P@�m���u�]��;]~��.���_^[��]� �����U���(W�}�����E�E���M��  �MS�؉EH����C�S�����E�ы���V�]�U��E܉U���]��~�E�E�K)}��]��'�M�U��E�Q�M�RP�����EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}�u�C�]��M���E�VP�҅��h����}�F���t)�M�+ȃ����    �Pf�\����f�f�u�]��}�;E�v����!���^[_��]� ��������U���(W�}�����E�E���M��,  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��:�M�E��M��t�M�+ȋ\�p���m���4u�EH�E����   )}��u�;E���$    �؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}�u�C�]��M��E�VP�҅��O����}�F���t%�M�+ȃ����    �\�P������u�]��}�;E�z�������^[_��]� ������������U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   |O���E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t}O�}�G�}��E9E�~�_^3�[��]� ��~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �������������U��V�u�F��F�����������������]�E�l  �]�����E��������D�Ez��^�P�P�]��������]��E����������N�X�N^�X]�����������U�������P�P��P�P�P�P �P�P�P,�P(�P$�U�M��U��U��U����M��U�P�ɋU��U��U��P�U�H�U��U��M����U��H�M��ɉP�U�U��]��H�M��P�U��]��P$�U��H �M��H(�P,��]�������������U���`�M�A,V�I�A(�I ���I�A(�I�A�I,���I���A�I �A�I���I$���]���E��������Dz�u�؋��������^��]���W���]�A�I,�A�I(�A�I�A�I �A(�I �U��A,�I�]������I$�����I�����e��	���E�������]��A�I�U��A�I�]��A�I,�]��A(�I�U����e��I$�E�������������A�������������]��A�I�A�I �����	�����A�������E��e��I���E�ʍu��ɋ��]��E��e����]��E��e����]����������]��A$�I �A�I,�����]��A,�I�A$�I�����]��A�I�A �I�����]��A(�I�A$�I�����]��A$�I�A(�I�����]��A�I�A�I�   �����]��_^��]�����������U�������P�P��P�P�X�خ�@    �U��U��U��]�M��Ԯ��M��U��U��P�]�U�P�U��H�M��H�P��]����������U��y t�U��������Au���B�A������Au�B�Y�B�A������Au�B�Y��A������z��Y�B�A������z�B�Y�B�A������z6�B�Y]� �E��Q�P�Q�@�A�Q�A��Q�A�Q�A   ]� ��������U����y ��   ��E�A�]��A�A�]��A�A�]��E��8������]�U��E�����]�U�P�M��]��U��P�A� �]��A�`�]�U��A�M��`�E��P�]��M��H��]� ��E�U�V�u��U�U��]�M��P�p�E��P�p^��]� �������������̋�3ɉ�H�H�H�V����t	P��<�����F�    ��t	P�<�����F    �F    �F    ^��U��V��W��t	P�}<�����F�    ��t	P�g<�����}�F    �F    �F    ����   �? ��   �G����   3ɺ   ����h�jlh�=���Q�~=�������t@� tB�G��t;3ɺ   ����h�jqh�=���Q�F=�����F��u�������_3�^]� �G��F�G��    Q�F�RP辠���F����t�N�W��QPR袠����_�   ^]� ����U��SV��W3�;�t	P�Z;�����F�>;�t	P�H;�����~�~�~9}�  �];��   3ɋú   ����h�h�   h�=���Q�q<�������tD9}tM�}��tF3ɋǺ   ����h�h�   h�=���Q�5<�����F��u�������_^3�[]� �~�73ɸ   �F�   ����h�h�   h�=���Q��;�����F��t���U��    PQR�^�x����E����t!�N�V��QRP�\�����_^�   []� �F�_^�   []� ������������3���A�A�A���U��Q�A�`�
�@�b�	���B�a����]��E���]�������U���|��UV�U��q�<��M��E�    �,  S�]W���  ��Uԋ�UЋM�U̍@�<����}��x�@�E��B�@�����E��}����>��U����]��@�E��������]��@�E��E��E؋E�����E����]ȋEȉE�   ;��  �w����`  �w�����F�B��   �U�P��R�������]��B���]��B�U����]��E����E������E��M������]��E��E������E����������]��E��M؉U؋U����ɉU܋U�U���P��R���]��E��E��]��E��E��]��E��E��]�����]��B���]��B���]��E����E������E��M������]��E��E������E��ˋU��������]��E��M؉U؋U����ɉU܋U�U����R���]��E��E��]��E��E��]��E��E��]�����]��B���]��B�U����]��E����E������E��M������]��E��E������E����������]��E��M؉U؋U����ɉU܋U�U��P��R���]��E��E��]��E��E��]��E��E��]���������]��B���]��B�U����]��E����E������E��M������]��E��E������E����������]��E��M؉U؋U����ɉU܋U�U����]��E��E��]��E��E��]��E��E��]��������U�E��;���   �ۍ�+���@����������]��@���]��@�E����]��E����E������E��M������]��E��E������E����������]��E��M؉E؋E����ɉE܋E�E����]��E��E��]��E��E��]��E��E��]��g�������������������UȋE��UċU��]��M���S�M�Q�U�R�C��������ẺK$�ыP�S(�@�C,������z	�����]��U�E�������z	�����]���U��E�E������E�����   ��������z���]��������z	�����]���U��E�E�������zb�������C(�����C,���]��M��C$���C,�����]ċU��c$�K�S�]ȋEȉC�C�K(�C�K,���]��C�K,�C�K$�   �����������z���]��������z���]��E�E���������   �C,�����C(���]��M��C$�����]ċU��C$���C(�K�ʉS���]ȋEȉC�C(�K�C,�K���]��C,�K�C$�K�M����]ċU��C$�K�C(�K�K�S���]ȋEȉC �{�C(�����C,�������]��M��K$�C,���]ċU��c(�K�S�]ȋEȉC �C�K,�C �K(���]��M��C$�K �C,�K���]ċU��C(�K�C$�K�K�S���]ȋEȉC�M�SQ������U�   �����M������3�3�3���|'�y�����B�U�҉U�U�w����u�U�};�}�Q���U��U�9��E�Ƌu�E����@�����K��@�K���@�K$���]��C��C�@�K���C(�H���]��C��C�@�K ���C,�H�E��E��E����E��]ȋEȉE��E��D��@�����K��@�K���@�K$���]�� �K�C�@�K���C(�H���]�� �K�C�@�K ���C,�H�ẺE����]ԋEЋI���EċE�3��Eȅ���   �F���FU�;���@�E�����K�U���@�K���@�K$���]��C��C�@�K���C(�H���]��C��C�@�K ���@�E��K,���]��E����E������E��U��U��ʉU��E��U����E���E��E��E��E��ʉU��ʉE��������E������]�E�E��]��5����E�_[^��]� �������h�=Ph_� �������������������h�=jh_� �o�������uË@����U��V�u�> t/h�=jh_� �C�������t��U�M�@R�Ѓ��    ^]���U��Vh�=jh_� ���	�������t�@��t�MQ����^]� 3�^]� �������U��Vh�=jh_� �����������t�@��t�MQ����^]� 3�^]� �������U��Vh�=jh_� ����������t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�=jh_� ���9�������t�@��t�MQ����^]� 3�^]� �������U��Vh�=j h_� �����������t�@ ��t�MQ����^]� 3�^]� �������U��Vh�=j$h_� ����������t�@$��t�MQ����^]� 2�^]� �������Vh�=j(h_� ���|�������t�@(��t��^��3�^������Vh�=j,h_� ���L�������t�@,��t��^��3�^������U��Vh�=j0h_� ����������t�@0��t�MQ����^]� 3�^]� �������U��Vh�=j4h_� �����������t�@4��t�M�UQR����^]� ���^]� ��Vh�=j8h_� ����������t�@8��t��^��3�^������U��Vh�=j<h_� ���i�������t�@<��t�MQ����^]� ��������������U��Vh�=j@h_� ���)�������t�@@��t�MQ����^]� ��������������U��Vh�=jDh_� �����������t�@D��t�MQ����^]� 3�^]� �������U��Vh�=jHh_� ����������t�@H��t�MQ����^]� ��������������Vh�=jLh_� ���l�������t�@L��t��^��3�^������Vh�=jPh_� ���<�������t�@P��t��^��^��������Vh�=jTh_� ����������t�@T��t��^��^��������Vh�=jXh_� �����������t�@X��t��^��^��������U��Vh�=j\h_� ����������t�@\��t�M�UQR����^]� 3�^]� ���U��Vh�=j`h_� ���i�������t�@`��t�M�UQR����^]� 3�^]� ���U��Vh�=jdh_� ���)�������t�@d��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh�=jhh_� �����������t�@h��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�=jlh_� ����������t�@l��t�M�UQR����^]� 3�^]� ���U��Vh�=jph_� ���I�������t�@p��t�M�UQR����^]� 3�^]� ���U��Vh�=jth_� ���	�������t�@t��t�M�UQR����^]� 3�^]� ���U��Vh�=jxh_� �����������t�@x��t�MQ����^]� 3�^]� �������U��Vh�=j|h_� ����������t�@|��t�M�UQR����^]� 3�^]� ���U��Vh�=h�   h_� ���F�������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�=h�   h_� �����������t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�=h�   h_� ����������t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���X��A�U�V�U��]����z  S��E��EW����������O  ���������U�r�z�
�R;��4v���I�$��4����R����   �]��F�a�]��F�a�]���!�]��B�a�]��B�a�]��E����E������E����E����������]��E������E������������]��������]��E��E��]��E��E��]��E��   �]��F�a�]��F�a����]���!�]��B�a�]��B�a�]��E����E������E����E����������]��E������E������������]��������]��E��E��]��E��E��]��E��E��]����m������_[�u�E�PV�|�������^��]� U���$V��M������F����   �6S�]W�u��E���$    ���������t[��%�����E�M܋���@��P�����F�@��R�M������~���Q�M��}����v;�t�v��P�M��g����u����m��u�u�_[�M�UQR�M�����^��]� ��������������̋Q3���|�	��t��~�    t@����u��3���������U��QV�u;��}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��|+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~#V�1�d$ ���   @u	�����t@����u�^���̋QV3���~�	�d$ ����ШtF����u��^���������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%���;��E���}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$���E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ���������������U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V����t	P�#�����F�    ��t	P�#�����F    �F    �F    ^��U��3�V���F�F�F�EP�������^]� �������������U��EVP��������^]� ����������U��SV��W3�;�t	P�#�����F�>;�t	P�#�����]�~�~�~;�tw3ɋú   ����h�jIh�=���Q�A$�������tJ�}��tL3ɋǺ   ����h�jNh�=���Q�$�����F��u���t	P�"�����    _^3�[]� �~_�^^�   []� ���U��Q�A�E� ��~LS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U�����u�_^[�E��Ћ�]� ���������U��3�V��W�}��F�F�F�Gj;Gu2j������tY�����O�H�G��B�N_���   ^]� j�f�����t'�����W�Q��O�H��G�B�N�   _��^]� ��̡�=�H��   ��U�존=�H��  V�u�R�Ѓ��    ^]����������̡�=�P��  Q�Ѓ�������������U�존=�P�EPQ��  �у�]� ̡�=�H�������U�존=�H�AV�u�R�Ѓ��    ^]��������������U�존=�H�AV�u�R�Ѓ��    ^]��������������U�존=�P��Vh�  Q���   �E�P�ы�=���   �Q8P�ҋ�=���   ��U�R�Ѓ���^��]��������������̡�=�P�BQ�Ѓ����������������U�존=�P�EPQ���   �у�]� �U�존=�P�EP�EP�EP�EP�EPQ���   �у�]� �U�존=�P�EP�EP�EP�EPQ�Jx�у�]� �������̡�=�P�B$Q��Y�U�존=�P�EP�EP�EP�EPQ��(  �у�]� �����U�존=�P�EP�EP�EPQ�J �у�]� ������������U�존=�H��8  ]��������������U�존=�P�EP�EP�EP�EPQ�J(�у�]� ��������U�존=�P�EP�EPQ�J,�у�]� U�존=�P�EP�EP�EPQ�J0�у�]� ������������U�존=�P�EP�EP�EP�EPQ�J<�у�]� ��������U�존=�P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U�존=�P�EP�EP�EP�EPQ�J@�у�]� ��������U�존=V��H�QWV�ҋ���=�H�QV�ҋ�=�Q�M�RHQ�MQ�MQOWHPj j V�҃�(_^]� ���������������U�존=�P�E P�EP�EP�EP�EP�EP�EPQ�JH�у� ]� ������������U�존=�P�EP�EPQ�JX�у�]� U�존=�P�EPQ�J\�у�]� ���̡�=�P�BlQ�Ѓ���������������̡�=�P�BlQ�Ѓ���������������̡�=�P�BpQ�Ѓ����������������U�존=�P�EPQ�Jt�у�]� ����U�존=�P�EPQ�Jt�у�]� ����U�존=�P�EP�EPQ���   �у�]� �������������U�존=�P�E���   ��VP�EPQ�M�Q�ҋu�    �F    ��=���   j P�BV�Ћ�=���   �
�E�P�у� ��^��]� ������̡�=�P���   Q�Ѓ���������������3��Yl��A`�Ad�Ah�Ap�����At   ����������������U��E��t�Al��yd t�Ah]� 3��yt��]� ������̡�=�H�������U�존=�H�AV�u�R�Ѓ��    ^]��������������U�존=�P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U�존=�P�EPQ�J�у�]� ���̡�=�P�BQ��Y�U�존=�P�EP�EPQ�J�у�]� U��VW�������M�U�x@�EPQR���n����H ���_^]� �U��VW���T����M�U�xD�EPQR���>����H ���_^]� �V���(����xH u3�^�W�������΍xH�����H �_^�����U��V��������xL u3�^]� W��������M�U�xL�EPQR��������H ���_^]� �������������U��V�������xP u3�^]� W�������M�U�xP�EP�EQRP���v����H ���_^]� ���������U��V���U����xT u3�^]� W���@����M�xT�EPQ���.����H ���_^]� �U���S�]VW���t.�M��&w����������xL�E�P��������H ��ҍM��w���}��tZ��=�H�A`�U�R�Ћ�=�Q�Jp�E�WP�ы�=�B�Pl�M�Q�҃��������@@��t��=�QWP�Bp�Ѓ�_^[��]� ������U��VW���d����xH�EP���V����H ���_^]� ���������U��VW���4����M�U�xD�EP�EQRP�������H ���_^]� �������������U��V��������xP u
�����^]� W��������M�U�xP�EP�EQ�MR�UPQR�������H ���_^]� ��������������U��V�������xT u
�����^]� W���}����M�xT�EPQ���k����H ���_^]� ��������������U��V���E����xX tW���7����xX�EP���)����H ���_^]� ������������U����MV3��E�PQ�u�u��u��u�u��  ����t.�E�;�t'��=�J�U�R�U�R�U�R�U�RP�Ax�Ѓ�^��]�3�^��]����������������VW���w���������3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_l��G`�Gd�Gh�Gp�����Gt   ��_^��������������V��W�>��t7�������xP t$S������j j �XPj�FP��������H ���[�    �~` t��=�H�V`�AR�Ѓ��F`    _^������������U��SV��Fp��=�Q��8  WV�^dSP�EP�~`W�у��Ft����   �> t�; ��   �U�~lW�^hSR�XC������u��h8�h�   ����I�����E�~P���+����j j jW�}����Ft��t��������Ft_^[]� �Ft_�Fp����^[]� �Ft�����    ��=�Q��JP�у��    �Ft_^[]� ��V��������3��^l��F`�Fd�Fh�Fp�����Ft   ^�������U��V��~d �F`t?W�};~pt5WPj�NQ�������Ft��u�F`�~p_^]� �M�Fp������t�3�_^]� �������������U��QVW�}����>  ��=�H���   V�҃���uh8�h�  �H����_3�^��]� ��=�E    �H�U�R�U�EP��  RV�Ѓ���t�3�9u�~"�E��I �<� t��Q���  �EF;u�|�UR������_�   ^��]� �������������U��QVW�}����~  ��=�H���   V�҃���uh8�h�  ��G����_3�^��]� ��=�E    �H�U�R�U�EP��  RV�Ѓ���tˋE��t�3�9u�~;��E�<� t*����=�QP���   �Ѓ���t�M��R���,  F;u�|ǍEP�����_�   ^��]� �������������h8�h�   h�=jx��������t�������3�����������V���8����N^�_������������������U��VW�}�7��t�������N�3���V������    _^]�h�=Ph�f � ������������������U��h�=jh�f ���������t
�@��t]�����]�������U��Vh�=jh�f ����������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�Z����E�NP�у�4�M���t�����^]ÍM�g������^]��U��h�=jh�f �<�������t
�@��t]��3�]��������U��h�=jh�f ��������t�x t�P]��3�]������V��FW��u�~��N�<��u�< ��u_3�^á�=�H�F���  h��j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� }(�V;Vu��������t�F�N��    �F9~|؋V;Vu���������t��F�N�U���F_�   ^]� ��������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T����H;ǉ�F�M���F_�   ^]� ����U��E��|2�Q;�}+J;Q}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�C��3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�د�M	��3����_�F�F^��������������U���SV�uW���^S�}��	��3���F�F�O�N�W���V9G�E~|��I �O���F�U�9FuL��u�~��~��t���< ��tY��=�H����  h��j8��    RP�у���t0�~�}���V��M����E�F@;G�E|�_^�   [��]� _^3�[��]� U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|���P�����_^]� �U����E�Qj�E��ARP�M��E���k�����]� �����U����Q�Ej�E��A�MRPQ�M��E��������]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q�����t!�A��t�B�A�Q�P�A    �A    �̋�� ��@���HV3��q�q�P�r�r����p�p�p�P�H^������V���������F3��F��;�t�N;�t�H�F�N�H�V�V�F�F��;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3����;�t�F;�t�A�F�N�H�V�V�Et	V��������^]� ������������U��V��W�~W�د���3����E��F�Ft	V�����_��^]� ������U��V��������Et	V�y������^]� ��U���V�u��u�a>  �@�E��0>  ���E�F�}� �E�u�E�H�����   �� ��   S�]W�   ;�s��uS�8  Y��u�   �F�Xt}��u�]��}��~7  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPW�u�j ��6  ��$��u������E�t	�M����_[^�Ë�U��V�^=  �@�u��+=  jh   �F�=  YY�F��th   �6  P�v��,  ���F   ��6  �f �F��^]Ë�Wh&������uV� >V��  ����`>Y|�^��_�h&����}V� >V�  ����`>Y|�^Ë�U��E��V��}k� >P�  Y��^]� ���}k� >P�  YË�U���u��0  Y��t]�<>  ]ËI������t�j���Ë�U��V��������EtV�!��Y��^]� ��U��E���t覥����t�j���]Ë�U��Qj �M��@���hh>������%h> Y�M��N����áh>Ë�U��=�> uhH���>��  Y�E�h>]�j�4��>  j �M�������}�e� �w��GN���8 t�������t�j�����w��w�  �M��Y�M��������>  Ë�U��Qj �M�������ȋ j�d>������d>��u�M������Ë�U��=d> uh�����Yj����Y��t�d>��M�H�3��d>]Ë�U��E�xP v�xTr�@@���@Pj �L  YY]�j�W��=  ��u��F   3��E��F�F�F�Eh���N���F�.������=  � j����o=  ��u���V�E�   ����Yj j�N�����H��=  Ë�U��V�������EtV���Y��^]� j����=  �h>����u{P�M��2����h>!u�����uXj4����Y�ȉM��E���t
V�������3�V�E� ������N�F?   �$����%���Ή5l>�����l>��>�M���M����������<  Ë�U��E�xVWr�p��pj j �!K  YY��u����}P�O<�%����tVj ��J  YY��u���P�OX�x%��_^]Ë�U��VW���w ��vW�u�V�6����u�_^]� ��U��V�uWj ��������F��t�8P���Y�ǅ�u�F �f ��t�8P���Y�ǅ�u�f  _^]Ë�U��V�u�~ v�F���>�F���> V����Y�N$��tj�y���^]Ë�Vj���J ��P��2  YY��^Ë�V���6�0  �6�)��YY^��1�.  Y��1�5  YË�U���V�u��u�8  �@�E���7  ���E�F�}� �E�u�E�H�����   �� ��   S�]��   s!��uS�@2  Y��u�   �F�X��   ��u�]��}�� 1  �M��H% �  ��N�]��}��E�%�   �A������t�E�j�E�]�E X�
3��]�E @j�u��M�jQP�EPh   �u�j �q0  ��$��u������E�t	�M����[^�Ë�U��V�u���(������^]� ���)����U��V�����)���EtV� ��Y��^]� jD�Ց��9  h��M���*���e� �E�P�M��(��h8��E�P��  �jD�Ց�9  h��M��*���e� �E�P�M��P���h�E�P�  ̋�U��V�u����1������^]� ��U��USVW�ڋ�����   ��@t����t��3Ɂ�;���3�A;�t��<�@��u�������8� u3��^��t%��t �uh4��u�	I  ����t	P�_  Y���u��h&V�u��H  ������t���tjj V��  ����tV�ŋ�_^[]Ë�U���  �'3ŉE��Eh  Ph  ������Pj �L  ����t3���u�������uP��������M�3���  �Ë�U���u� �]Ë�U���u�$�]Ë�U���u�(�]Ë�U���u�,�]Ë�U�졬&��u]�6  �MH��&���>]�����>@��&��t���>��&��
r������̋L$WSV��|$��to�q��tU���L$���:�t��t���:�t
��u�^[_3�Ê��:�u�~��a��t(���:�u��A��t�f���:�t��3�^[_���K  �G�^[_Ë�^[_Ë�U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$����U��QQSVWd�5    �u��E���j �u�u��u�J} �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u��V  �� �E�_^[�E���]Ë�U��V��u�N3��  j V�v�vj �u�v�u�V  �� ^]Ë�U���8S�}#  u����M�3�@�   �e� �E���'�M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E��Y  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M�  �E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u�eU  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����-���u�9\  �M�N��k���M9H};H~���u	�M�]�u�} }ʋEF�0�E�;_w;�v��[  ��k�E�_^[�Ë�U��EV�u��DX  ���   �F�6X  ���   ��^]Ë�U���!X  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V��W  �u;��   u��W  �N���   ^]���W  ���   �	�H;�t���x u�^]�J[  �N�H�ҋ�U����'�e� �M�3��M�E��E�E�E@�E�	��M��E�d�    �E�E�d�    �uQ�u�C[  �ȋE�d�    ����;'u���q[  ��Q�Ȱ�i\  YË�U��V��������EtV�����Y��^]� ��U��E��	Q��	P�\  ��Y�Y@]� ��U��E��t���8��  uP�J  Y]Ë�U��EV���F ��uc�V  �F�Hl��Hh�N�;.t�0-�Hpu��5  ��F;8,t�F�0-�Hpu��^  �F�F�@pu�Hp�F�
���@�F��^]� ��U����'3ŉE�S3�V;�u�c  j^SSSSS�0�  ���5  �uW�)c  YY;Er��ЋU��H;�u ��8t�<a|<z, �A8u�3���   j�p�   SSj�WVQR��'  �ȃ�$�M�;�u�)c  � *   �c  � �   9Ms��c  j"�^���;�~Ej�3�X���r9�A=   w�;c  ��;�t� ��  �P�a  Y;�t	� ��  ���M�E���]�9]�u�b  �    냋U�j�pQ�u�j�WV�pR� '  ��$��t�u��uW��   ������lb  j*Y����u������Y�ƍe�^[�M�3��}����Ë�U���W�u�M�������}�E�P�u�_����}� YY_t�M��ap��Ë�U��j �u�u������]Ë�U��S3�9D?uA�E;�u��a  SSSSS�    �H	  ��3��/��8t)�
��a|
��z�� �
B8u��Sj��u�X����E��[]Ë�U��MS3�VW;�t�};�w�{a  j^�0SSSSS��  �����0�u;�u��ڋъ�BF:�tOu�;�u��@a  j"Y�����3�_^[]������̋T$�L$��ti3��D$��u��   r�=D[ t��a  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�ø�g��/��/�^��/t^��/�^��/^��/��/Qg��/2^��/�]��/!]Ë�U��������m  �} � ?t�Sm  ��]���U��WV�u�M�}�����;�v;���  ��   r�=D[ tWV����;�^_u^_]�n  ��   u������r*��$�D���Ǻ   ��r����$�X��$�T���$����h�����#ъ��F�G�F���G������r���$�D��I #ъ��F���G������r���$�D��#ъ���������r���$�D��I ;�(� ���� ����D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�D���T�\�h�|��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$����I �Ǻ   ��r��+��$����$�������@��F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I �����������������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë��` �` � ܰË�U��S�]VW���ܰ���t&P�;)  ��FV�  YY�G��t�3VP���������g �G   ��_^[]� ��U��S�]V���ܰ�C�F���CWt1��t'P��(  ��GW�  YY�F��t�sWP�������	�f ��F_��^[]� �y �ܰt	�q��  YËA��u��Ë�U��V�EP�����������^]� ��U��V�u���R��������^]� ���������U��V�������EtV�����Y��^]� ��U��V������c����EtV����Y��^]� ��U��V�uW3�;�u3��e9}u�5[  j^�0WWWWW�  �����E9}t9urV�u�u�/  �����uW�u�������9}t�9us��Z  j"Y����jX_^]������������̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[Ë�U��EVW3�;�tG9}u�Z  j^�0WWWWW�k  �����)9}t�9Es��Y  j"Y�����P�u�u������3�_^]Ë�U��E�$?]Ë�U���(  �'3ŉE������� SjL������j P�Z�����������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   �������D�j ���@���(���P�<���u��uj��g  Yh ��8�P�4��M�3�[�����Ë�U���5$?�H  Y��t]��j�g  Y]����3�PPPPP�������Ë�U��� �EVWjY���}��E��E_�E�^��t� t�E� @��E�P�u��u��u��H��� jhH�9t  �u��tu�=<[uCj�+i  Y�e� V�Si  Y�E��t	VP�ti  YY�E������   �}� u7�u�
j�h  Y�Vj �5�B�P���u�W  ���L�P�@W  �Y��s  �jhh�s  3��}�3��u;���;�u �UW  �    WWWWW����������   V�=v  Y�}��F@uwV��z  Y���t���t�����ȃ���� J��p3�A$u)���t���t��������� J��p3�@$�t��V  �    WWWWW�1������M��9}�u�Nx
��A��V�v  Y�E��E������   �E��s  ËuV��u  Y�jh��r  3��}�3��u;���;�u �QV  �    WWWWW����������   V�9u  Y�}��F@uwV��y  Y���t���t�����ȃ���� J��p3�A$u)���t���t��������� J��p3�@$�t��U  �    WWWWW�-������M��9}�u!�Nx��E�����V�u�ty  YY�E��E������   �E���q  ËuV��t  YË�U��V�u�F@WuyV�y  Y�p3���t���t�ȃ�������� J����A$u&���t���t�ȃ������ J����@$�t��T  3�WWWWW�    �_���������JS�]���t=�F�u��y2�u.3�9~uV�z  Y�;Fu9~u@���F@�t8t@����[_^]È�F�F�����F��%�   ��jh��p  3�3�9u��;�u�YT  �    VVVVV�����������+�u�Bs  Y�u��u�u�����YY�E��E������	   �E��p  ��u�s  YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�w  YP葀  ��;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�w  P��  Y��Y��3�^]�jh��o  3��}�}�j�d  Y�}�3��u�;5 [��   � K��98t^� �@�tVPV�Ur  YY3�B�U�� K���H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u� K�4�V�^r  YY��E������   �}�E�t�E��	o  �j��b  Y�jh��n  3�9uu	V����Y�'�u�aq  Y�u��u����Y�E��E������	   �E��n  ��u�q  Y�j�����Y�jh	�Rn  3ۉ]�3��u;���;�u ��Q  �    SSSSS�c���������   �E��t	;�t��@u�;�t��@u�}�G�=���v뷋}����uV�p  Y�]�V����V��  YY�f�����N�Et���Fj_�-�E;�u W��  Y;�u�$D�M����N  �	��   �N�~�F��^�E������	   �E��m  ��u�p  YË�U���SVW3�9}t$9}t�u;�u��P  WWWWW�    �f�����3�_^[�ËM;�tڃ��3��u9Ew͋}�}�F  �M��}��t�F�E���E�   ����   �N��  t/�F��t(��   ��;�r��W�u��6�  )~>��+�}��O;]�rO��tV�S���Y��u}�}� ��t	3ҋ��u�+�W�u�V��s  YP��|  �����ta��;�w��M�+�;�rP�}��)�E�� VP��s  YY���t)�E��FK�E����E�   ���A����E������N ��+�3��u������N �E���jh0	��k  3�9ut)9ut$3�9u��;�u �O  �    VVVVV�������3�� l  ��u�}n  Y�u��u�u�u�u�=������E��E������   �E����u�n  YË�U��W3�9}u�,O  WWWWW�    ����������AV�u;�u�O  WWWWW�    �n����������u��  Y�ȉ#ʃ���V;�t3�^_]Ë�U��V�u�F��u�N  �    ����g���}�FuV�9�  E�e YV�����FY��y����F��t�t�   u�F   �u�uV�r  YP��  3Ƀ������I��^]�jhP	�xj  3�3�9u��;�u�'N  �    VVVVV����������>�};�t
��t��u��u��l  Y�u�W�u�u�������E��E������	   �E��Oj  ��u�?m  YË�U��V3�9uu�M  VVVVV�    �����������E;�t�V�p�0�u�V�  ��^]Ë�U��SV�uW3����;�u�cM  WWWWW�    ���������B�F�t7V�:���V���{  V��p  P��  ����}�����F;�t
P����Y�~�~��_^[]�jhp	�7i  �M��3��u3�;���;�u��L  �    WWWWW�G����������F@t�~�E��:i  �V�k  Y�}�V�*���Y�E��E������   �ՋuV�l  YË�U��Q�e� S�]��u3��   W��ru�{���vn�M�E�������tR:Q�uM�P���t<:Q�u7�P���t&:Q�u!�P���t:Q�u�E�9}�r��?�@��I��F�@��I��<�@��I��2�@��I��(�M�E����t:u@A�E�9]�r�3�_[��� �	+����U���u�T���u�L��3���tP��K  Y���]�3�]Ë�U��� WV�0  3�Y;�u�~K  WWWWW�    �����������49}t޹����E�I   �u�u��M�;�w�E��u�E��u�uP�U��_�Ë�U��V�u�EPj �uhP��z�����^]Ë�U��j
j �u�>�  ��]Ë�U��EVW��u|P�	Z  Y��u3��  �?  ��u�Z  ��諜  �\��H[�d�  �,?�k  ��}�;  ��菚  ��| ��  ��|j �ߕ  Y��u�(?�   ��m  ��3�;�u19=(?~��(?9=TDu�n�  9}u{�m  �#;  �Y  �j��uY��:  h  j��  ��YY;��6���V�5�'�5P?�9:  Y�Ѕ�tWV�;  YY�X��N���V�����Y�������uW�=  Y3�@_^]� jh�	��e  ����]3�@�E��u9(?��   �e� ;�t��u.�$���tWVS�ЉE�}� ��   WVS�r����E����   WVS�|����E��u$��u WPS�h���Wj S�B����$���tWj S�Ѕ�t��u&WVS�"�����u!E�}� t�$���tWVS�ЉE��E������E���E��	PQ�w�  YYËe��E�����3��Pe  Ë�U��}u�r�  �u�M�U�����Y]� ��������������̃=�I ���  ���\$�D$%�  =�  u�<$f�$f��f���d$�l�  � �~D$f(@�f(�f(�fs�4f~�fTp�f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�,�  ���D$��~D$f��f(�f��=�  |!=2  �fT0��\�f�L$�D$����f�`�fV`�fTP�f�\$�D$���������������̃=D[ t-U�������$�,$�Ã=D[ t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$��jh�	��b  �e� �u;5,[w"j��W  Y�e� V��_  Y�E��E������	   �E���b  �j��V  YË�U��V�u�����   SW�=`��=�B u�؟  j�&�  h�   �(�  YY�<[��u��t���3�@P���uV�S���Y��u��uF�����Vj �5�B�׋؅�u.j^9�Ht�u趟  Y��t�u�{�����E  �0��E  �0_��[�V菟  Y�E  �    3�^]Ë�U��� S3�9]u�E  SSSSS�    �����������N�E;�t�V�u�E��u�E��u�E�P�E�����E�B   ��  ���M��x�E����E�PS�i  YY��^[�Ë�U���uj �u�u�m�����]����̀�@s�� s����Ë����������������������������U��WV�u�M�}�����;�v;���  ��   r�=D[ tWV����;�^_u^_]��R  ��   u������r*��$����Ǻ   ��r����$���$����$�(���#ъ��F�G�F���G������r���$���I #ъ��F���G������r���$���#ъ���������r���$���I �xph`XPH�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�0�����$���I �Ǻ   ��r��+��$�4�$�0�Dh��F#шG��������r�����$�0�I �F#шG�F���G������r�����$�0��F#шG�F�G�F���G�������V�������$�0�I ����'�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�0��@HXl�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_���5�H�1  Y��t��j�A�  jj �  ���|  ��U��QSVW�5�I�o1  �5�I���}��_1  ��YY;���   ��+ߍC��rwW�ը  ���CY;�sH�   ;�s���;�rP�u���  YY��u�G;�r@P�u���  YY��t1��P�4��z0  Y��I�u�l0  ���V�a0  Y��I�EY�3�_^[�Ë�Vjj �=  ��V�:0  ����I��I��ujX^Ã& 3�^�jh�	�\  �X�  �e� �u�����Y�E��E������	   �E��\  ��7�  Ë�U���u���������YH]���̺`'��  �`'�l�  �Ƀ= ?t���贶  �����z�����������������̃��$���  �   ��ÍT$診  R��<$�D$tQf�<$t�`�  �   �u���=? �Ӻ  �   ��'�к  �  �u,��� u%�|$ u���5�  �"��� u�|$ u�%   �t����-�4�   �=? �v�  �   ��'��  ZË�U����'3ŉE�SV3�W��9<?u8SS3�GWh��h   S�p���t�=<?��L���xu
�<?   9]~"�M�EI8t@;�u�����E+�H;E}@�E�<?����  ;���  ����  �]�9] u��@�E �5l�3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�l>  ��;�t� ��  �P����Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �5p�SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�=  ��;�tj���  ���P�����Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�p���t"SS9]uSS��u�u�u�VS�u �h��E�V�z���Y�u��q����E�Y�Y  �]�]�9]u��@�E9] u��@�E �u��  Y�E���u3��!  ;E ��   SS�MQ�uP�u ��  ���E�;�tԋ5d�SS�uP�u�u�։E�;�u3��   ~=���w8��=   w�<  ��;�t����  ���P����Y;�t	� ��  �����3�;�t��u�SW��������u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��]�  ���u������#u�W�O���Y��u�u�u�u�u�u�d���9]�t	�u�����Y�E�;�t9EtP�y���Y�ƍe�_^[�M�3������Ë�U����u�M��
����u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap����-  �ȋAl;.t�0-�Qpu�  ���   Ë�U����u�M������E����   ~�E�Pj�u��  ������   �M�H���}� t�M��ap��Ë�U��=D? u�E�.�A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u萸  ������   �M�H���}� t�M��ap��Ë�U��=D? u�E�.�A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Pj�u��  ������   �M�H���}� t�M��ap��Ë�U��=D? u�E�.�A��]�j �u����YY]Ë�U����u�M������E����   ~�E�Ph�   �u菷  ������   �M�H%�   �}� t�M��ap��Ë�U��=D? u�E�.�A%�   ]�j �u�~���YY]Ë�U����u�M������E����   ~�E�Pj�u��  ������   �M�H���}� t�M��ap��Ë�U��=D? u�E�.�A��]�j �u����YY]Ë�U���L�'3ŉE�S3�V�uW�]ԉ]�]��]؉]܉u��]�9^�  �F9u P�F0h  P�E�SP�e�  ������  j�  j��  W�E��  jW�E��  jW�E��  jh  �E��  ��$�E�9]��|  9]��s  ;��k  9]��b  9]��Y  �Eԉ3��M܈@=   |�E�P�v�t����/  �}��%  �E���E�~-8]�t(�E�:�t�x�����M�� �G;�~�@@8X�uۋE�SS�v   Ph   �u܉E�jS�ѷ  �� ����  �M��E�S�v��   W���   QW@Ph   �vS������$����  �E�S�v�   WP�E�W@Ph   �vS�U�����$���`  �E�}����   3҃}�f��U؉Mč��   �_�Z��M����   �MȈ~S8]�tN�M�M�:�tB�I���;ʉM�'��H   ��M��E� �  f�AA�M̋M��	9M�~�M�AA�M�8Y�u�h�   ��   QP�=���j��   PW�.����E�j��   QP�������   ��$;�tKP����u@���   -�   P��������   ��   +�P�������   +�P�������   �������E��    ���   �E����   �Eĉ��   �E����   �Eȉ��   �EЉ��   �u��S���Y���m�u��F����u��>����u��6����u��.���3ۃ�C�ˍ��   �;�tP������   ǆ�   ��ǆ�   �ǆ�   ��ǆ�      3��M�_^3�[�������X'  �ȋAl;.t�0-�Qpu�r  �@��2'  �ȋAl;.t�0-�Qpu�L  ��Ë�U��VW3��u������Y��u'9@?vV�����  ;@?v��������uʋ�_^]Ë�U��VW3�j �u�u�%�  ������u'9@?vV�����  ;@?v��������uË�_^]Ë�U��VW3��u�u���  ��YY��u,9Et'9@?vV�����  ;@?v��������u���_^]Ë�U��VW3��u�u�u�÷  ������u,9Et'9@?vV�����  ;@?v��������u���_^]��̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+�Ë�U���(  �'3ŉE���'Vtj
莊  Y蟷  ��tj衷  Y��'��   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P���������������(�����0���j ǅ����  @��������,����@���(���P�<�j��~  ̋�U��M��'�U#U��#�ʉ�']�Pd�5    �D$+d$SVW�(��'3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(��'3�P�e��u��E������E�d�    ËM�d�    Y__^[��]QË�U��SV�u���   3�W;�to=�6th���   ;�t^9uZ���   ;�t9uP��������   ���  YY���   ;�t9uP�������   落  YY���   �������   ����YY���   ;�tD9u@���   -�   P�n������   ��   +�P�[������   +�P�M������   �B��������   �= 6t9��   uP���  �7����YY�~P�E   ��8-t�;�t9uP�����Y9_�t�G;�t9uP�����Y���Mu�V�����Y_^[]Ë�U��SV�5�W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�8-t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5�W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{�8-t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�V���t��t;�tWj6Y���  P����Y_^Å�t7��t3V�0;�t(W�8����Y��tV�����> Yu��@-tV�3���Y��^�3��jh�	�wJ  �   ��0-�Fpt"�~l t�   �pl��uj �x  Y���J  �j�F?  Y�e� �Fl�=.�i����E��E������   ��j�A>  Y�u�á.�H��B�H��B���   �.���   ��6���   �7���   ��'���   �7�3�Ë�U��SW�}3�;�~,V�u���6�u�u蚿  ����tSSSSS������Ou�^_[]Ë�U��SVW�}h�   3�SW������u�����u3���   <.u4�F8t-jP���   jP���  ����tSSSSS�/��������   ��h��V�]荿  ;��   �} �<0�u��@��   ��.��   PVj@�u�;�}u��@sw��_trP�EVj@��@��}u`��s[��t��,uRP�EVj��P�f�  ����t3�PPPPP��������,�'����������E�wh��V��  ��YY�X������_^[]Ë�U��SV�uV�u�u�b�����3ۅ�tSSSSS�6������F@8tPh��j�u�u�Q��������   8^[tPh��j�u�u�/�����]Ë�U���S3�ChU  �]������Y�E���U  W�x� ��]��^�CH�0�E�h���5ܹjhQ  W������E���E��E�ܹh��hQ  W�t�  ����t3�PPPPP�k������sX�E��0�B#  YY��t�e� �E��E��E����0�CH�0�E�E�h���0jhQ  W�Z������}��|��}� uI�FP����tP�Ӆ�u	�vP����Y�FT��tP�Ӆ�u	�vT����Y�E�fT �fL �FP�~H���N�u��i����FP�=�3�Y;�tP�ׅ�u	�vP�J���Y�FT;�tP�ׅ�u	�vT�3���Y�Fh�^T�^L�^P�^H_[�Ë�U���   �'3ŉE��ESV�uW�}��d����E��\�����`����o  �   �H(��T����H,�X �   ��X�����h�������  ��d��� ��  �} ��  �>CuW�~ uQh���u��d����������3���tVVVVV�������;�t3�f�f�Gf�G��`���;�t�0��d����G  V�������   Y��P���;�s,V��h����_!  YY����   V��X����I!  YY����   ��L��� ��l���VP����YY����   ��l���PSP�Y�  ������   �C��T������l���PW��h����������> t
��P���;�r��L������@PVW��X���蓻  ����t3�VVVVV��������3�9�\���tjS��\����}�����9�`���tj��T�����`����_�������h����u��d�����������tVVVVV�`�������h����3��M�_^3�[�)����Ë�U����  �'3ŉE�SW���[  �u����h���P��P���Ph�   ��x���PS���  ��������u3��  �E���0�sH��x���P�  YY���x  ��x���P������P��t��������YY��p�����t��CH�M��\����D���k���l���� ��X����1jP��d�����<���P�?����F��x���Q��t�����L�����p��������QP�X�������t3�PPPPP�,�������p�����l������CH��P����j��P���P��d�����������}��   ��h�����t��� �F�G$�O ��d����ǋV;t6���t������d�����D����P�H��D�������t�����d���|��"��t�����t�ǋ��P�W���d����H��t���uhj�v��x����vPjh�jj 誦  �� ��t93���  f!�Ex���@��r�h�   �5�'��x���P�3�  �����@�G��g �F��G���   �}u	��h����F�Ek�V��عY��t1��\�����p����CH�k�����X���Y��l������L����F������\���8-t-�E�����<0�7����u�7�#����sT�����cL YY�M��p��������    �1�CH�M�_3�[�'����Ë�U���   �'3ŉE��ESV3ۋ�W��h���;�t;�tP�����Y��  ���D0H��  ǅp���   ��t���;���  �9L�0  �yC�&  �y_�  ��h��W�b�  ��YY����   +ǉ�p�����   �;;��   ǅl���   �ܹ���p���PW�6��������u�6�����Y9�p���t��l��������~�Ch��S軶  ��3�YY;�u	�;;��   ��l���QWS��x���h�   P�Ҷ  ����tVVVVV��������l�����h�����x���Ƅ=x��� ����Y��t��t�����? t
G�? � ���3�9�t�����   ��h����u3��vSSSh�   ��x���PQ�"�����;�tZ�~H��t3�7��x���P�b  YY��tS��x����%���Y��u!�p������t���C����~�3�9�p���u9�t���t�D����M�_^3�[������jh
�
?  3ۉ]��}v�"  �    SSSSS�#�����3��,  �!  ���u��N����Np�]�jh�   �8���YY���}�;���   j�3  Y�E�   �Nl�������]��   �u�M���P���Y�E�;���   9]th8-�u�[  YY��t
�D?   j�U3  Y�E�   �^l���y���W����Y�Fpu2�0-u)�;�.�W���j�.��Ph�B�������������e� �   �-�}܋u�3�j�2  YËu�j�2  Y��W�K���W�m���YY�E������   �E���=  Ëu�fp��jhH
�=  3��u�3��];���;�u�D!  �    VVVVV������3��{3��};���;�t�3�f97��;�t����  �E;�u�!  �    �ɉu�f93u ��   �    j��E�Ph'���  ���P�uWS���  ���E��E������	   �E��0=  ��u� @  YË�U���SV�u3ۉ]�;�t9]u3��{  v3�f�W�};�u�l   SSSSS�    ��������<  �u�M�������E�;���   9XuH9]v�M��9f�f�8tAFF�M�;Mr�8]�t�E�`p��E���   8]�t�E�`p�����   �uVj�W�=l�j	�p��;���   �L���zt��  � *   3�f��   �E�u�E�;�t'��M�:�t�M���QP��  YY��tF8t!F9]�u��u+u�u�E�V�uj�p��;�uT�a  �M� *   3�f��-9Xu	W�����Y�1SSj�Wj	�p�l�;�u�*  � *   8]�t�E�`p�����H8]�t�M�ap�_^[�Ë�U���SV�u3ۉ]�;�u9]t*�9]w��  j^SSSSS�0�B���������   3�f�W�};�t��u�M��Y����E;Ev�E=���v	�  j�P�M�QP�uV����������u;�t3�f��h  � 8]�tk�M�ap��b@;�tH;Ev<�}�t,3�f��>  j"^SSSSS�0������8]�t�E�`p����&�E�E�P   3�f�LF�;�t�8]�t�E�`p��E�_^[�Ë�U��j �u�u�u�u�u�������]�������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[Ë�U��V�EP���7��������^]� ����������U��V����������EtV�����Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR�  YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =MOC�t=csm�u+�  ���    ��  �  ���    ~�  �   �3�]�jhh
�68  �}�]��   �s��s�u��\  �   � �e� ;ute���~;w|��  �����Oȋ1�u��E�   �y t�sh  S�O�t��  �e� ��u��-���YËe�e� �}�]�u��u���E������   ;ut�a  �s��7  Ë]�u��  ���    ~�  �   �Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�q  3�A��  ���3��jh�
�7  �M��t*�9csm�u"�A��t�@��t�e� P�q�&����E������7  �3�8E��Ëe��R  ̋�U��M�V�uƃy |�Q�I�42���^]Ë�U�����u
�c  �  �e� �? �E� ~SSV�E�@�@��p��~3�E����E�M�q�P�GE�P�_�������u
K�������E��E��E�;|�^[�E���j���u����X  ���    t��  �e� �  �M���|  �3  �Mj j ���   �J����j,h��5  �ً}�u�]�e� �G��E��v�E�P蜳��YY�E���  ���   �E���  ���   �E���  ���   ��  �M���   �e� 3�@�E�E��u�uS�uW�������E�e� �o�E������Ëe��  ��   �u�}�~�   �O��O�^�e� �E�;Fsk�ËP;�~@;H;�F�L�QVj W�������e� �e� �u�E������E    �   �E��5  ��E�맋}�u�E܉G��u�����Y��
  �Mԉ��   ��
  �MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v�j���Y��t�uV�%���YY�jh0�24  3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w�b�  YY����   SV�Q�  YY����   �G��M��QP�����YY���   �}�E�p�tH��  YY����   SV�	�  YY����   �w�E�pV���������   ���t|��W�9Wu8���  YY��taSV���  YY��tT�w��W�E�p�_���YYPV赶�����9��  YY��t)SV��  YY��t�w�z�  Y��t�j X��@�E���  �E������E��3�@Ëe��Q  3��3  �jhP�2  �E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS衭����FP�w����YYP�vS臭���E������2  �3�@Ëe��  ̋�U��} t�uSV�u�V������}  �uuV��u �E����7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP�Ϭ��]Ë�U��QQV�u�>  ���   W��  ���    t?��  ���   �z  9t+�>MOC�t#�u$�u �u�u�u�uV�i���������   �}� u�"  �u�E�P�E�PV�u W豮�����E���;E�s[S;7|G;wB�G�O����H��t�y u*�X��@u"�u$�u�u j �u�u�u�u�����u���E��E���;E�r�[_^�Ë�U���,�MS�]�C=�   VW�E� �I��I����M�|;�|�h
  �u�csm�9>��  �~� ��  �F;�t=!�t="���   �~ ��   �  ���    ��  �  ���   �u�q  ���   jV�E��  YY��u��	  9>u&�~u �F;�t=!�t="�u�~ u�	  �&  ���    t|�  ���   �  �u3����   ����Y��uO3�9~�G�Lh�'�Ϯ����uF��;7|��	  j�u�d���YYh���M��7���hl�E�P�Һ���u�csm�9>��  �~�~  �F;�t=!�t="��e  �}� ��   �E�P�E�P�u��u W艬�������E�;E���   �E�9��   ;G|�G�E�G�E��~l�F�@�X� �E��~#�v�P�u�E����������u�M��9E���M�E��}� ��(�u$�]��u �E��u��u�u�uV�u�K����u���E����]����}�} t
jV�:���YY�}� ��   �%���=!���   �����   V����Y����   �_  �Z  �U  ���   �J  �}$ �M���   Vu�u��u$�.����uj�V�u�u�������v�����]�{ v&�} �)����u$�u �u�S�u�u�uV������� ��  ���    t�_  _^[�Ë�U��V�u���մ�������^]� ��U��SVW�  ��   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������� 3�@_^[]Ë�U��V�5�'�5���օ�t!��'���tP�5�'���Ѕ�t���  �'�ܺV�x���uV�aZ  Y��th̺P�|���t�u�ЉE�E^]�j ����YË�U��V�5�'�5���օ�t!��'���tP�5�'���Ѕ�t���  �'�ܺV�x���uV��Y  Y��th��P�|���t�u�ЉE�E^]����� ��V�5�'�������u�5L?�e���Y��V�5�'�����^á�'���tP�5T?�;���Y�Ѓ�'���'���tP�����'���  jh��+  �ܺV�x���uV�'Y  Y�E�u�F\��3�G�~��t$h̺P�|��Ӊ��  h���u��Ӊ��  �~pƆ�   CƆK  C�Fh(j�  Y�e� �vh���E������>   j�  Y�}��E�Fl��u�.�Fl�vl�O���Y�E������   �*  �3�G�uj�m  Y�j�d  YË�VW�L��5�'�������Ћ���uNh  j������YY��t:V�5�'�5P?�����Y�Ѕ�tj V�����YY�X��N���	V脵��Y3�W���_��^Ë�V��������uj�X  Y��^�jh��)  �u����   �F$��tP�7���Y�F,��tP�)���Y�F4��tP����Y�F<��tP����Y�F@��tP�����Y�FD��tP����Y�FH��tP����Y�F\=��tP�Ҵ��Yj�  Y�e� �~h��tW����u��(tW襴��Y�E������W   j��  Y�E�   �~l��t#W�A���Y;=.t��@-t�? uW�M���Y�E������   V�M���Y��(  � �uj�  YËuj�  YË�U��=�'�tK�} u'V�5�'�5���օ�t�5�'�5�'���ЉE^j �5�'�5P?����Y���u�x�����'���t	j P���]Ë�VW�ܺV�x���uV�V  Y�����^  �5|�h(�W��h�W�H?��h�W�L?��h�W�P?�փ=H? �5���T?t�=L? t�=P? t��u$����L?����H?�K�5P?�T?�����'�����   �5L?P�օ���   �%X  �5H?�����5L?�H?�����5P?�L?�����5T?�P?�u������T?�v  ��teh�M�5H?�����Y�У�'���tHh  j�6�����YY��t4V�5�'�5P?����Y�Ѕ�tj V�y���YY�X��N��3�@��$���3�_^�jh��j&  �����@x��t�e� ���3�@Ëe��E������6����&  ��~����@|��t������jh�&  �5X?����Y��t�e� ���3�@Ëe��E������}����h�P�g���Y�X?����������U���SQ�E���E��EU�u�M�m��U�  VW��_^��]�MU���   u�   Q�3�  ]Y[�� ��U���(  �h@�d@�`@�\@�5X@�=T@f��@f�t@f�P@f�L@f�%H@f�-D@��x@�E �l@�E�p@�E�|@��������?  �p@�l?�`?	 ��d?   �'�������'�������D���?j�  Yj �@�h4��<��=�? uj�|  Yh	 ��8�P�4���jh8�z$  j�|  Y�e� �u�N��t/��B��B�E��t9u,�H�JP�����Y�v�����Y�f �E������
   �i$  Ë���j�G  Y��������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�ҥ��3��ȋ��~�~�~����~����(���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �'3ŉE�SW������P�v�t��   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R������C�C��u�j �v�������vPW������Pjj 迆  3�S�v������WPW������PW�vS������DS�v������WPW������Ph   �vS�^�����$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[�P�����jhX�N!  �������0-�Gpt�l t�wh��uj �O  Y���f!  �j�"  Y�e� �wh�u�;58,t6��tV����u��(tV褬��Y�8,�Gh�58,�u�V���E������   뎋u�j��  YË�U���S3�S�M�������B���u��B   ���8]�tE�M��ap��<���u��B   ����ۃ��u�E��@��B   ��8]�t�E��`p���[�Ë�U��� �'3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�@,��   �E��0=�   r����  �p  ����  �d  ��P������R  �E�PW�t����3  h  �CVP�/���3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�����M��k�0�u���P,�u��*�F��t(�>����E���<,D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C��D,Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95�B�X�������M�_^3�[�K�����jhx�I  �M���������}�������_h�u�u����E;C�W  h   �J���Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh����u�Fh=(tP耩��Y�^hS�=����Fp��   �0-��   j�  Y�e� �C��B�C��B�C��B3��E��}f�LCf�E�B@��3��E�=  }�L��0*@��3��E�=   }��  ��8+@���58,����u�8,=(tP�Ǩ��Y�8,S���E������   �0j�  Y��%���u ��(tS葨��Y�   �    ��e� �E��  Ã=�I uj��V���Y��I   3�Ë�U��3�9Ev�M�9 t@A;Er�]Ë�U��E3�;�(.tA��-r�H��wjX]Ë�,.]�D���jY;��#���]�������u��/Ã���������u��/Ã�Ë�U��V������MQ�����Y�������0^]��������������Q�L$+ȃ����Y骸  Q�L$+ȃ����Y锸  U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh���  �e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E���  Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[�������D[3�Ë�U���V�u�M��w����u�P�A�  ��e�F�P�������Yu��P�$�  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�`�  �M��E��M��H��EP��  �E�M����Ë�U��j �u�u�u������]Ë�V����tV����@PV�V�(�����^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M��������3�;�u+����j_VVVVV�8�l������}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�����j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h<�SV詙����3ۅ�tSSSSS�}������N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F��Ht�90uj�APQ襚�����}� t�E��`p�3�_^[�Ë�U���,�'3ŉE��ESVW�}j^V�M�Q�M�Q�p�0��  3ۃ�;�u�y���SSSSS�0���������o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q��  ��;�t���u�E�SP�u��V�u��������M�_^3�[�����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �U���9}}�}�u;�u+����j^WWWWW�0��������}� t�E�`p����  9}vЋE��� 9Ew	�Q���j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV��  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� �Ͷ  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �y�  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V������u�E�8 u���} �4����$�p���WF��  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP��  0�F�U�����;�u��|��drj jdRP躴  0��U�F����;�u��|��
rj j
RP蔴  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N������u-�.���j^�03�PPPPP蔝�����}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V�K������}� t�E��`p�3�_^[�Ë�U���,�'3ŉE��ESVW�}j^V�M�Q�M�Q�p�0譲  3ۃ�;�u����SSSSS�0芜�������Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P�ְ  ��;�t���u�E�SV�u���`������M�_^3�[�׏���Ë�U���0�'3ŉE��ESV�uWj_W�M�Q�M�Q�p�0��  3ۃ�;�u�d���SSSSS�8�ϛ�������   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW��  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[�ݎ���Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3����/�6������Y���(r�_^Ë�Vh   h   3�V��  ����tVVVVV������^Ë�U����P��]��H��]��E��u��M��m��]����]�����z3�@��3���ht������thX�P�|���tj �������U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]Ã%@[ Ë�U��3�9Ej ��h   P�����B��u]�3�@�<[]Ã=<[uWS3�9$[W�=P�~3V�5([��h �  j �v�����6j �5�B�׃�C;$[|�^�5([j �5�B��_[�5�B����%�B Ë�VW3���B�<��/u���/�8h�  �0��衯  YY��tF��$|�3�@_^Ã$��/ 3����S�$�V��/W�>��t�~tW��W辗���& Y�����0|ܾ�/_���t	�~uP�Ӄ����0|�^[Ë�U��E�4��/�,�]�jh��  3�G�}�3�9�Bu��H  j�9G  h�   �;:  YY�u�4��/9t���nj袺��Y��;�u�#����    3��Qj
�Y   Y�]�9u,h�  W蘮  YY��uW����Y������    �]���>�W�і��Y�E������	   �E��F  �j
�(���YË�U��EV�4��/�> uP�"���Y��uj�/9  Y�6�(�^]Ë�U��$[�([k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   � D����   �8[�5��h @  ��H� �  SQ�֋8[� D�   ���	P� D�@�8[����    � D�@�HC� D�H�yC u	�`�� D�x�ueSj �p�֡ D�pj �5�B�P��$[� Dk��([+ȍL�Q�HQP�K����E���$[; Dv�m�([�0[�E� D�=8[[_^�á4[V�5$[W3�;�u4��k�P�5([W�5�B���;�u3��x�4[�5$[�([k�5([h�A  j�5�B�`��F;�t�jh    h   W����F;�u�vW�5�B�P�뛃N��>�~�$[�F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�����u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U����$[�Mk�([������M���SI�� VW}�����M���������3���U��0[����S�;#U�#��u
���];�r�;�u�([��S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1�([�	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t�0[�C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u; Du�M�;8[u�% D �M���B_^[��h�wd�5    �D$�l$�l$+�SVW�'1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q���������������̋�U���S�]V�s35'W��E� �E�   �{���t�N�38�S~���N�F�38�C~���E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t�����  �E���|@G�E��؃��u΀}� t$����t�N�38��}���N�V�3:��}���E�_^[��]��E�    �ɋM�9csm�u)�=�� t h����  ����t�UjR������M胙  �E9Xth'W�Ӌ�膙  �E�M��H����t�N�38�=}���N�V�3:�-}���E��H����  �����9S�R���h'W���1�  ������0á [Vj^��u�   �;�}�ƣ [jP�Y���YY� K��ujV�5 [�@���YY� K��ujX^�3ҹ�0�� K��� ����p3|�j�^3ҹ 1W������ J����������t;�t��u�1�� B��`1|�_3�^������=PD t�W�  �5 K����YË�U��V�u��0;�r"��P3w��+�����Q�����N �  Y�
�� V�(�^]Ë�U��E��}��P������E�H �  Y]ËE�� P�(�]Ë�U��E��0;�r=P3w�`���+�����P�����Y]Ã� P�,�]Ë�U��M���E}�`�����Q����Y]Ã� P�,�]Ë�U��V�uW3�;�u����WWWWW�    �k�������   �F����   �@��   �t�� �F��   ���F�  u	V�  Y��F��v�vV�W  YP�P�  ���F;���   �����   �F�uOV�-  Y���t.V�!  Y���t"V�  ��V�<� J�  ��Y��Y��p3�@$�<�u�N    �~   u�F�t�   u�F   ��N�A���������	F�~���_^]�jTh�� ���3��}��E�P�Ġ�E�����j@j ^V�y���YY;��  � J�5�I��   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@� J��   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M��� J���I ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=�I|���=�I�e� ��~m�E����tV���tQ��tK�uQ�����t<�u���������4� J�E� ���Fh�  �FP��  YY����   �F�E�C�E�9}�|�3ۋ���5 J����t���t�N��r�F���uj�X�
��H������P��������tC��t?W�����t4�>%�   ��u�N@�	��u�Nh�  �FP�y�  YY��t7�F�
�N@�����C���g����5�I���3��3�@Ëe��E������������Ë�VW� J�>��t1��   �� t
�GP�$����@   ;�r��6�W����& Y���� K|�_^Ë�U��EV3�;�u�8���VVVVV�    蟃���������@^]Ë�U��QV�uV�����E�FY��u������ 	   �N ����/  �@t������ "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,������� ;�t�������@;�u�u�Х  Y��uV��   Y�F  W��   �F�>�H��N+�I;��N~WP�u�  ���E��M�� �F����y�M���t���t����������� J��p3�@ tjSSQ�1�  #����t%�F�M��3�GW�EP�u�  ���E�9}�t	�N �����E%�   _[^�Ë�U���$Dh   ����Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U���  �t�  �'3ŉE��EV3���4�����8�����0���9uu3���  ;�u'�:����0� ���VVVVV�    臁��������  SW�}�����4� J�����ǊX$�����(�����'�����t��u0�M����u&�����3��0����VVVVV�    �������C  �@ tjj j �u�:�  ���u�ͣ  Y����  ��D���  ������@l3�9H�������P��4�� ����Р���`  3�9� ���t���P  �̠��4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P�^�  Y��t:��4���+�M3�@;���  j��@���SP��  �������  C��D����jS��@���P��  �������  3�PPj�M�Qj��@���QP�����C��D����h������\  j ��<���PV�E�P��(���� �4�Ƞ���)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4�Ƞ����  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@������  Yf;�@����h  ��8����� ��� t)jXP��@����ҡ  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4�Ƞ���B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4�Ƞ���b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �h���;���   j ��,���P��+�P��5����P��(���� �4�Ƞ��t�,���;����L���@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0�Ƞ��t��,�����@��� ��8�����L���@�����8��� ul��@��� t-j^9�@���u����� 	   �����0�?��@�������Y�1��(�����D@t��4����8u3��$�h����    �p����  ������8���+�0���_[�M�3�^�nn����jh��l����E���u�4����  ����� 	   ����   3�;�|;�Ir!�����8������ 	   WWWWW�Xz�����ɋ����� J��������L1��t�P�ݠ  Y�}���D0t�u�u�u�.������E������� 	   �����8�M���E������	   �E��������u�'�  Y�jh�����E���u�E���� 	   ����   3�;�|;�Ir�$���� 	   SSSSS�y�����Ћ����<� J��������L��t�P��  Y�]���Dt1�u脟  YP�Ԡ��u�L��E���]�9]�t������M������ 	   �M���E������	   �E�������u�F�  YË�U��V�u�F��t�t�v�Zy���f����3�Y��F�F^]Ë�U��   �S�  �'3ŉE�SV�uWV�������3�9FY������}�FjPPS�@�  ������������������|��s
������  ������ J��������� ��ÊH$����F  ������u�F�������+�ʋǋ��  ��V��+��V���������Z  �������  3�9P0�  �����9Vu�������������<  R�p,�p(�������o�  ��������� Ã���;p(�0���;x,�'���j ������Qh   ������Q�0�ؠ������j ��������������������  ����������������������������;��������������t7������K;�s+���u�J�;�s�H�9
u�������07�@��uЍ�����+�3����L  �@�t�V��:
u������B;�r������������u�������  ��x������    �$����F��   �V��u!�������   +N��@�����   jj j ��������  ��;�����u$;�����u�F�8��8
uG@;�r��F    �Yj �������������������×  �����������������   ;�w�N��t
����   t�~������� �DtG������u��)����������� ������uѭ����������3������������M�_^3�[�4i����jh8�2����u�����Y�e� �u����Y�E��U��E������   �E��U��D�����u�4���YË�U��V�uV�W�  Y���u����� 	   ����MW�uj �uP�ܠ�����u�L��3���tP����Y���������� J�����D0� ���_^]�jhX�s����E���u�;����  � ���� 	   ����   3�;�|;�Ir!�����8������ 	   WWWWW�_t�����ɋ����� J��������L1��t�P��  Y�}���D0t�u�u�u��������E������� 	   �����8�M���E������	   �E��������u�.�  YË�U���SW�}3�;�u �M���SSSSS�    �s��������f  W�����9_Y�E�}�_jSP�������;ÉE�|ӋW��  u+G�.  ��OV��+�u���tA�U��u����� J�����D2�t��;�s���:
u�E�3�B;�r�9]�u�E���   ��x������    �   �G��   �W;�u�]��   �]��u�+�������� J�E����D0�tyjj �u�������;E�u �G�M��	�8
u�E@;�r��G    �@j �u��u����������}����:�   9Ew�O��t��   t�G�E��D0t�E�E)E��E�M��^_[�Ë�U��V�u�FW��ty�}��t
��t��uh���F��uV�I���EYU3�V�v���FY��y����F��t�t�   u�F   W�u�uV����YP肓  #����t3���9����    ���_^]�jhx�^����u�!���Y�e� �u�u�u�u�:������E��E������	   �E��k�����u�[���YË�U��V�uWV�}�  Y���tP� J��u	���   u��u�@Dtj�R�  j���I�  YY;�tV�=�  YP� ���u
�L����3�V虖  ������ J����Y�D0 ��tW�s���Y����3�_^]�jh��s����E���u�;����  � ���� 	   ����   3�;�|;�Ir!�����8������ 	   WWWWW�_p�����ɋ����� J��������L1��t�P��  Y�}���D0t�u�����Y�E������� 	   �M���E������	   �E�������u�=�  YË�U��9EuF�jP;Mu+����YY���u3�]ËE�    �6�u�7�^������Q��������tՉ�&3�@]Ë�U���EP�`������EYu��߃�]��Jx	�
�A�
�R�����YË�U��}�t]�mr��]Ë�U��S�U�������؃��t��P����Y��u��[]Ë�U����  �'3ŉE��M�EV3�W�}�������|�����d�����T���ǅ$���^  ��0����������x���;�u �K���VVVVV�    �n��������5  ;�t��@@SuzP�����Y�p3���t���t�ȃ�������� J����A$u&���t���t�ȃ������ J����@$�t �����VVVVV�    �-n��������  �u������Ob���ƅc��� ��t�����<������k  ��d�����P�ȍ��Y��t0��t���VV��t�������YP�k���YYG�P蝍��Y��u��  �<%�1  8G�  3���@���ƅ/��� ��X�����L�����l���ƅa��� ƅ`��� ƅj��� ƅS��� ƅb��� ƅs��� ƅk�����(���G���P����Y��t��l�����L���k�
�DЉ�l�����   ��N��   ��   ��*tp��F��   ��It��Lut��k����   �O��6u�G�84u��(�������4�����8����m��3u�G�82u���\��dtW��itR��otM��xtH��Xu�A��j����9��ht(��lt��wt��S����"�G�8lt���k�����s������k�����s�����S��� �������j��� ��H���u������0�������������3�2ۉ�D���8�s���u�<Stƅs����<Cuƅs������ ��\�����ntJ��ct��{t��d�����t����}���Y���d�����t����@�����x��������  ��D�����H�����L�����t��l��� ��  ��\�����o�r  �  ��c�
  jdZ;���  �z  ��g~E��it!��n�g  ��j��� ��t����f
  �
  ��\�����x���-�4  ƅ`����1  3ۃ�x���-u��T���� -C�	��x���+u��l�����d�����t����^�����x�����L��� u��l������x����k��l�����l�����tf��x�����T�����X������0���P��|���PCS��T�����$�������������
  ��d�����t����������x�����P����Y��u���������   � � ��a���:�x�����   ��l�����l�������   ��d�����t���������T�����x�����a������0���P��|���PCS��T�����$��������������	  ��x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$����{���������	  ��d�����t����������x�����P����Y��u���X��� �_  ��x���et��x���E�I  ��l�����l������5  ��T����e��0���P��|���PCS��T�����$��������������  ��d�����t����D�����x�����-u,��T����-��0���P��|���PCS����������  �	��x���+u/��l�����l�����u!�l������d�����t����������x�����x����k��l�����l�����tf��T�����x�����X������0���P��|���PCS��T�����$������������  ��d�����t����j�����x�����P誆��Y��u���d�����t�����x����U�����X��� YY��  ��j��� ��  ��T�����<��������QP��D���� ��k���HP�5�/�&���Y�Ѓ��  ��u��l���ǅL���   ��s��� ~ƅb�����d�����t���W��x�����@�������YY��L��� t��l�����l������3  ��t������x�����x�������  ��\���ctN��\���su��	|	����  �� u2��\���{��  ��a���3ҋȃ�B������L�3˅���  ��j��� ��  ��b��� �~  �� �����P�v  Y��t��t������������!��������P�����ǅ���?   ���   �� ���P�����P��  f�������f�FF�  ��p��  �������HH�{  ���������t3�;�x�����  ��c�����j��� �  �����������  ��s��� ~ƅb���G�?^��u
�wƅa����j �E�j P��\�����>]u	�]F�E� �f��/����^F<-uB��t>���]t7F:�s�����:�w"*������Ћσ��ǳ�����D�GJu�2���ȊЋ��������D��<]u����  ��H�����D���������x���+u'��l���u��t����d�����t����C�����x���j0^9�x����x  ��d�����t���������x���<xtX<XtT��\���xǅX���   t"��L��� t
��l���u��ǅ\���o   �$  ��d�����t���P�����YY��x����  ��d�����t���������L��� ��x���t��l�����l���}��ǅ\���x   ��   �F��D����������@���������t���WP�j���YY9�@�����  ��j��� �  ��<�����\���c��  ��b��� t��D���3�f���  ��D����  ��  ƅk�����x���-u	ƅ`����	��x���+u'��l���u��t����d�����t���������x�����(��� �J  ���  ��\���xte��\���pt\��x���P�с��Y����   ��\���ou"��x���8��   ��4�����8��������Rj j
��8�����4����̋  �����7��x���P�����Y��tr��4�����8�����x������������Y��x�����x�����X�����Й����L��� ��4�����8���t��l���t5��d�����t���������x���������d�����t�����x�������YY��`��� ��@�����   ��4�����8����؃� �ى�4�����8�����   ��@�������   ��\���xt;��\���pt2��x���P聀��Y����   ��\���ou��x���8}n���,k�
�'��x���P�Ӏ��Y��tR��x����������Y��x�����X�����L��� ��x����|�t��l���t5��d�����t���������x����X�����d�����t�����x�������YY��`��� t�߃�\���Fu��X��� ��X��� �  ��j��� u8��<�����D�����(��� t��4������8����F���k��� t�>�f�>��H�����c���G��H����`<%u
�G�8%u����t�������������G��x�����H���;�ul��P�p  Y��t!��t�����������G��H���;�uG��t�����x����u�?%uD��H����xnu8������	����*��d�����x�������YY�VS��VP����VS�y�������0���u��T����B`��Y��x����u*��<�����u8�c���u�������� t%������ap������� t
������`p���<���[�M�_3�^�!S���Ë�U���VW�u�M��S���E�u3�;�t�0;�u,�����WWWWW�    �(_�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�5  �M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&� ����E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9D?uh .�P������]Ë�U��W��  W���u�x����  ��`�  w��t�_]Ë�U����  �u�6  �5�3�~���h�   �Ѓ�]Ë�U��h���x���th��P�|���t�u��]Ë�U���u�����Y�u���j�7���Y�j�T���YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=̰ th̰�"u  Y��t
�u�̰Y�z���h��hx�����YY��uBh
��5t���\��$t��c����=�I Yth�I��t  Y��tj jj ��I3�]�jh��Q���j�S���Y�e� 3�C9XD��   �TD�E�PD�} ��   �5�I����Y���}؅�tx�5�I�����Y���u܉}�u����u�;�rW�ԣ��9t�;�rJ�6�Σ����辣������5�I踣�����5�I諣����9}�u9E�t�}�}؉E����u܋}��h������_���Yh������O���Y�E������   �} u(�XDj����Y�u�����3�C�} tj�h���Y��w���Ë�U��j j�u�������]�jj j ������Ë�V�������V�  V�Br  V��X��V�i  V��  V�G7  V��Q��V����h��G�����$��3^Ã=�I u�����V�5,?W3���u����   <=tGV��~��Y�t���u�jGW��}����YY�=8D��tˋ5,?S�BV��~����C�>=Yt1jS��}��YY���tNVSP�gP������t3�PPPPP�;X�������> u��5,?��Y���%,? �' ��I   3�Y[_^��58D�Y���%8D ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF��  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�0�  Y��t��M�E�F��M��E����  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9�Iu�q���h  �`DVS�dE���H[�5HD;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P��z����Y;�t)�U��E�P�WV�}�������E���H�,D�50D3�����_^[�Ë�U��hE��SV�5��W3�3�;�u.�֋�;�t�hE   �#�L���xu
jX�hE��hE����   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5h�SSS+�S��@PWSS�E��։E�;�t/P�z��Y�E�;�t!SS�u�P�u�WSS�օ�u�u��V��Y�]��]�W�����\��t;�u�����;��r���8t
@8u�@8u�+�@P�E��y����Y;�uV���E����u�VW�Mi����V����_^[�Ë�V������W��;�s���t�Ѓ�;�r�_^Ë�V������W��;�s���t�Ѓ�;�r�_^Ë�U��QQV�ȟ�������F  �V\��3W�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ��3�=�3���;�}$k��~\�d9 �=�3��3B߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]Ë�U����'�e� �e� SW�N�@��  ��;�t��t	�У'�`V�E�P���u�3u�� �3��X�3����3��E�P����E�3E�3�;�u�O�@����u������5'�։5'^_[�Ë�U���(3�S�]V�uW�}�E��E��E��E��E��E��E��E�9lEt�5�I諛��Y��~-�M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �E�ܼ��M��]�Q��]���]���Y����  ����� "   �  �E�ؼ��M��]�Q��E�   �]���]���Y�j  �E�   �E�ؼ��E�м��]���]���"  �M��E�м�r����E�̼�׉M��E�̼�Z����E�ܼ놃�tNIt?It0It ��t����   �E�ļ��Eܼ���E�ܼ����E�ܼ�x����E�   ��������   �E�   �Eܴ���������������   �$�±�E�̼��E�м��E�ؼ��Eܬ���Eܤ���Eܜ��y����Eܔ��m����Eܐ���E܌���E܈���M����]���]�M��]�Q�E�   ��Y��u�H���� !   �E��_^[��)�2�;�D�M�V��b�˰°n�w����%�I 谪����I3�Ë�U��QQSV���  V�5�3�5�  �EYY�M�ظ�  #�QQ�$f;�uU�ہ  YY��~-��~��u#�ESQQ�$j�]�  ���rVS��  �EYY�d�ES�`����\$�E�$jj�?�F�  �]��EY�]�Y����DzVS观  �E�YY�"�� u��E�S���\$�E�$jj�>�  ��^[�Ë�U��QQS�]VW3�3��}�;��3t	G�}���r���w  j蠄  Y���4  j菄  Y��u�=8?�  ���   �A  h���  S�pEW�F������tVVVVV��M����h  ��EVj ��F ����u&hp�h�  V��E������t3�PPPPP�M����V��s��@Y��<v8V��s����;�j��Hhl�+�QP�':  ����t3�VVVVV�WM�����3�hh�SW�:9  ����tVVVVV�3M�����E��4��3SW�9  ����tVVVVV�M����h  h@�W���  ���2j������;�t$���tj �E�P�4��3�6�&s��YP�6S�Ƞ_^[��j�$�  Y��tj��  Y��u�=8?uh�   �)���h�   ����YYË�U��E��H]Ë�U���5�H�P���Y��t�u��Y��t3�@]�3�]��A@t�y t$�Ix��������QP�����YY���u	��Ë�U��V����M�E�M�����>�t�} �^]Ë�U���G@SV����t2� u,�E�+��M���}���C�>�u�r����8*u�ϰ?�d����} �^[]Ë�U���x  �'3ŉE�S�]V�u3�W�}�u�������������������������������������������������������������@����u5�����    3�PPPPP�OL���������� t
�������`p������
  �F@u^V�b���Y�p3���t���t�ȃ�������� J����A$u����t���t�ȃ������ J����@$��g���3�;��]�������������������������������
  C������ �������
  ��, <Xw��������3��3�3������j��Y������;���	  �$����������������������������������������������v	  �� tJ��t6��t%HHt���W	  �������K	  �������?	  �������3	  �������   �$	  �������	  ��*u,����������;���������  ��������������  ������k�
�ʍDЉ�������  ��������  ��*u&����������;���������  ��������  ������k�
�ʍDЉ������{  ��ItU��htD��lt��w�c  ������   �T  �;luC������   �������9  �������-  ������ �!  �<6u�{4uCC������ �  ��������  <3u�{2uCC�����������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������P��P�������6Y  Y��������Yt"�����������������C������������������������������M  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@9������������   �������������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  ����������������  ;�u��4������������ǅ����   �  ��X��  HHty+��'���HH��  ��������  ������t0�G�Ph   ������P������P�~  ����tǅ����   ��G�������ǅ����   �������������5  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  ��4������P�5l��Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�7���������,|  ���/��������� tf������f���������ǅ����   �  ������@ǅ����
   �������� �  ��  ��W����  u��gueǅ����   �Y9�����~�������������   ~?��������]  V��i��������Y��������t���������������
ǅ�����   3�����������G�������������P��������������������P������������SP�5�/�D���Y�Ћ���������   t 9�����u������PS�5�/����Y��YY������gu;�u������PS�5�/�����Y��YY�;-u������   C������S����ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �i���������Qƅ����0������ǅ����   �E�����   �K������� t��������@t�G���G����G���@t��3҉�������@t;�|;�s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�'m  ��0��9����������~������N뽍E�+�F������   ������������ta��t�΀90tV�������������0@�>If90t@@;�u�+��������(;�u��4�������������I�8 t@;�u�+����������������� �\  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+�����������u������������Sj �p������������������������������v���������Yt������uWSj0�������.����������� ������tf��~b�������������������Pj�E�P������FPF�Cy  ����u(9�����t �������������M������������ Yu����������������P�����������Y������ |������tWSj ������������������ t�������1B�������� Y���������������t������������������������� t
�������`p��������M�_^3�[�5���Ð#�$�T�����	�O�}���U���   �'3ŉE��ESV�u3ۃ}W��t�����l�����   Sh�   ��|�����Q�u��x����uP�y  ����;�uj�L���z��   SSS�u�u��t����Wy  ����p���;�t_3�FVP��d����YY;�tMS��p�����x���W�u�u��t����y  ����;�tjV�d��YY��l����;�u!9�x���tW��@��Y����M�_^3�[��3���ÍN�QWVP��+  ����tSSSSS��>����9�x���tW�@��Y3��9]u�Sj��HW�u�uP�w  ����t�����P�^��Y��tɊ�
���,0GG���H�|�뱋�U��E��H]�jh��f���3��]3�;���;�u�����    WWWWW�z?��������S�=<[u8j�2���Y�}�S�[���Y�E�;�t�s���	�u���u��E������%   9}�uSW�5�B�������&����3��]�u�j� ���Y��������U���0���S�ٽ\�����=@8 t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=@8 t�#  ��8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq����,  �   [�À�8�����=? uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �8������������(�����s4�H��,ǅr���   �0������������ �����v�@�VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P��u  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����D   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Àzuf��\���������?�f�?f��^���٭^�����4�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����4�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����4���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-�4��p��� ƅp���
��
�t����������l$�l$�D$���   5   �   t��������4 u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t��4����4���l$�����4����4���l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r ��������4�|$�l$�ɛ�l$������l$��Ã�,��?�$�5����,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  �������4 �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����5�Ƀ�u�\$0�|$(���l$�-5�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8��4�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w����4�|$��4�<$� �|$$�D$$   �D$(�l$(����4�<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  �������4 �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u�����5�Ƀ�u�\$0�|$(���l$�-5�����l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8��4�l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w����4�|$��4�<$� �|$$�D$$   �D$(�l$(����4�<$�l$$�Q�����0Z�����0Z�������@���������������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�e  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   ��P��   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��|������������l������   s������t������������d������   v����떋�U����'3ŉE�j�E�Ph  �u�E� ����u����
�E�P�u8��Y�M�3�����Ë�U���4�'3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5t��M�QP�֋l���t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u��O����YF;�~[�����wS�D6=   w/�$�����;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�.<��Y;�t	� ��  ���E���}�9}�t؍6PW�u��L!����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�h���t`�]��[�h�9}�uWWWWV�u�W�u�Ӌ�;�t<Vj��M��YY�E�;�t+WWVPV�u�W�u��;�u�u���)��Y�}���}��t�MЉ�u��i��Y�E��e�_^[�M�3������Ë�U���S�u�M��_���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P��8  YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP��  �� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U��QQ�'3ŉE���HSV3�W��;�u:�E�P3�FVh��V����t�5�H�4�L���xu
jX��H���H����   ;���   ����   �]�9]u��@�E�5l�3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w蓀����;�t� ��  �P�9��Y;�t	� ��  ���؅�ti�?Pj S������WS�u�uj�u�օ�t�uPS�u���E�S�n���E�Y�u3�9]u��@�E9]u��@�E�u�����Y���u3��G;EtSS�MQ�uP�u��������;�t܉u�u�u�u�u�u����;�tV�]'��Y�Ǎe�_^[�M�3�����Ë�U����u�M������u$�M��u �u�u�u�u�u�������}� t�M��ap���jh��?����M3�;�v.j�X3���;E�@u��~���    WWWWW�K&����3���   �M��u;�u3�F3ۉ]���wi�=<[uK������u�E;,[w7j�ӏ��Y�}��u�ٗ��Y�E��E������_   �]�;�t�uWS�5����;�uaVj�5�B�`���;�uL9=�Ht3V����Y���r����E;��P����    �E���3��uj�w���Y�;�u�E;�t�    ���s����jh�!����]��u�u�d7��Y��  �u��uS�%��Y�  �=<[��  3��}�����  j�����Y�}�S�	���Y�E�;���   ;5,[wIVSP��������t�]��5V躖��Y�E�;�t'�C�H;�r��PS�u��k8��S蹎���E�SP�ߎ����9}�uH;�u3�F�u������uVW�5�B�`��E�;�t �C�H;�r��PS�u��8��S�u�蒎�����E������.   �}� u1��uF������uVSj �5�B�������u�]j����YË}����   9=�Ht,V�a���Y��������{|��9}�ul���L�P�&|��Y��_����   �V|��9}�th�    �q��uFVSj �5�B�������uV9�Ht4V�����Y��t���v�V�����Y�
|���    3�耘�����{���|�����u��{�����L�P�{���Y���ҋ�U��MS3�;�v(j�3�X��;Es�{��SSSSS�    �#����3��A�MVW��9]t�u�T���Y��V�u������YY��t;�s+�Vj �S�9������_^[]Ë�U��E��H��H��H��H]Ë�U��E��3V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5�H�1k��Y�j h8�)���3��}�}؋]��Lt��jY+�t"+�t+�td+�uD��l�����}؅�u����a  ��H��H�`�w\���]���������Z�Ã�t<��t+Ht�{z���    3�PPPPP��!����뮾�H��H���H��H�
��H��H�E�   P�mj���E�Y3��}���   9E�uj�&���9E�tP�U���Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.��3�M܋�3��3�9M�}�M�k��W\�D�E�����i����E������   ��u�wdS�U�Y��]�}؃}� tj ����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3��˕��Ë�U����HB�PD�M��U���u����Ãe� SW�E��FPj1Q3�C�E�SP�I������FPj2�u��E�SP�4�����FPj3�u��E�SP������FPj4�u��E�SP�
�����P��FPj5�u��E�SP�������FPj6�u��E�SP�����Vj7�u���E�SP�������F Pj*�u��E�SP������P��F$Pj+�u��E�SP������F(Pj,�u��E�SP������F,Pj-�u��E�SP�t�����F0Pj.�u��E�SP�_�����P��F4Pj/�u��E�SP�G�����FPj0�u��E�SP�2�����F8PjD�u��E�SP������F<PjE�u��E�SP������P��F@PjF�u��E�SP�������FDPjG�u��E�SP�������FHPjH�u��E�SP�������FLPjI�u��E�SP������P��FPPjJ�u��E�SP������FTPjK�u��E�SP������FXPjL�u��E�SP�o�����F\PjM�u��E�SP�Z�����P��F`PjN�u��E�SP�B�����FdPjO�u��E�SP�-�����FhPj8�u��E�SP������FlPj9�u��E�SP������P��FpPj:�u��E�SP�������FtPj;�u��E�SP�������FxPj<�u��E�SP�������F|Pj=�u��E�SP������P����   Pj>�u��E�SP��������   Pj?�u��E�SP�y�������   Pj@�u�S�E�P�a�������   PjA�u��E�SP�I�����P����   PjB�u��E�SP�.�������   PjC�u��E�SP��������   Pj(�u��E�SP���������   Pj)�u��E�SP�������P����   Pj�u��E�SP���������   Pj �u��E�SP��������   Ph  �u��E�SP��������   Ph	  �]�S�E�j P�{�����P���_���   [�Ë�U��V�u����  �v����v����v�����v�����v�����v�����6�����v �����v$�����v(�����v,����v0����v4����v����v8����v<�����@�v@����vD����vH�z���vL�r���vP�j���vT�b���vX�Z���v\�R���v`�J���vd�B���vh�:���vl�2���vp�*���vt�"���vx����v|�����@���   ������   �������   �������   �������   �������   �������   �������   ������   ������   ������   �����,^]Ë�U��SVW�}�  � 6t@h�   j�-?����YY��u3�@�E��������tV�+���V�J��YY��ǆ�      �����   �;�t�   P���73�_^[]Ë�U��V�u��t5�;�6tP����Y�F;�6tP����Y�v;5�6tV����Y^]Ë�U���S�]V3�W�]�u�9su9su�u��u��E�6�:  j0j�V>����YY�};�u3�@�w  ���   jYj���=��3�Y�E�;�u�u�`��Y�щ09s��   j��=��Y�E�;�u3�F�u�8���u��0��YY���  �0�u�{>VjW�E�jP�T����E�FPjW�E�jP�?���	E�FPjW�E��E�jP�'�����<E�tV����Y���뎋E�� ����0|��9��0�@�8 u��7��;u���~�����> u����6�E���6�H��6�u��H�E�3�A��E���t����   �5���tP�֋��   ��tP�օ�u���   �7�����   �,��YY�E����   �E����   �E���   3�_^[�Ë�U��V�u��t~�F;�6tP����Y�F;�6tP����Y�F;�6tP����Y�F;�6tP���Y�F;�6tP���Y�F ; 7tP���Y�v$;57tV�~��Y^]Ë�U���SV�uW3��}��u��}�9~u9~u�}��}���6�6  j0j��;����YY;�u3�@�u  j�;��Y�E�;�u	S���Y���89~��  j�~;��Y�E�;�uS�����u�����Y�҉8�v8�CPjV�E�jP�������CPjV�E�jP������CPjV�E�jP�������CPjV�E�jP�������P��CPjV�E�jP�������C PjPV�E�jP������C$PjQV�E�jP������C(PjV�E�j P������P��C)PjVj �E�P�r�����C*PjTV�E�j P�^�����C+PjUV�E�j P�J�����C,PjVV�E�j P�6�����P��C-PjWV�E�j P������C.PjRV�E�j P������C/PjSV�E�j P�������<�t$S����S����u�����u�������Q����C����0|��9��0�@�8 u��#��;u���~�����> u���jY��6���E�u�   ��	���I�K� �@�M��C3�@3��9}�t�M�����   ;�tP�����   ;�t#P����u���   �������   ����YY�E����   �E����   ���   3�_^[�Ë�U��ES3�VW;�t�};�w�m��j^�0SSSSS��������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u��Wm��j"Y����3�_^[]��������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^�Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w��l��j^�0SSSSS�*��������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x�����Hl��j"Y���낋�U��3�S3�@9]|FVW��t>�EÙ+��E���<��7�E�0�N  YY��u
�M���9�}N�u��^;]~�_^3Ʌ���[��]Ë�U����'3ŉE�V���tS�> tNh��V��c��YY��t=h��V��c��YY��uj�E�Pj�w����t/�u�V�r ��Y�M�3�^�����j�E�Ph  �w����u3��׍E�h��P�}c��YY��u����뻋�U��3�f�Mf;���t@@��r�3�@]�3�]Ë�V3��#��,aB<w������,A<w��������tЊ
��u׋�^�3��
B��A|��Z~��a��w@��Ë�U���|�'3ŉE�VW�}�.]�����ׁƜ   ������jx�E�P�F���%���  PW����u!F@�2�E�P�v�M  YY��uW����Y��t
�N�~�~�F���Ѓ��M�_3�^�d���� ��U���|�'3ŉE�Vjx�E�P�E%�  j   P������u3��.�U������9Et�} t�6W�������V���v6��Y;�_t�3�@�M�3�^�����Ë�U���|�'3ŉE�SVW�}�!\�����ׁƜ   �y�������jx�E�P�F���%���  PW�Ӆ�u�f 3�@�b  �E�P�v��K  YY����   jx�E�P�F���%���  PW�Ӆ�t��E�P�6�K  YY��u�N  �~�R�FuO�F��t,P�E�P�6��L  ����u�6�N�~�5��Y;Fu!�~��V��uW����Y��t	���V�~�N�   #�;���   jx�E�P�F���%���  PW�Ӆ������E�P�6�K  Y3�Y��u/�N   �F9^t
   �F�G9^t;�6��4��Y;Fu.j�9^u49^t/�E�P�6��J  YY��uSW�������YY��t�N   9^u�~�F���Ѓ��M�_^3�[����� ��U���|�'3ŉE�VW�}�PZ�����ׁƜ   ������jx�E�P�F���%���  PW����u!F@�[�E�P�6�)J  YY��u	9Fu0j��~ u0�~ t*�E�P�6�J  YY��uPW���$���YY��t
�N�~�~�F���Ѓ��M�_3�^�]���� �6��3���v�����@�F�3��������f @�~ YY�FtjX���	���jh@��F���F�   t�   t�u�f ��6�_3�������@Y�FtjX������jh��F���Fu�f Ë�U��SVW��X���]���Ɯ   ��u�N  �   �C@�~����t�8 tWjh�����������f ��tS�8 tN���t�8 t�������S����~ ��   Vj@h����������tb�?��t�? t�����P�����I�?��t0�? t+W�q2������Y�j@h4��F���Fu�f ��F  ���F�F�~ ��   �˃����#ˋ��������}����   ����  ��   ����  ��   ��P�������   j�v� �����   �E��tf�Nf�f�Nf�Hf�x�]��tm�=��  f9u%h��j@S�W������t"3�PPPPP�+�����j@Sh  �v�ׅ�t,j@�C@Ph  �v�ׅ�tj
j��S�u��I  ��3�@�3�_^[]Ë�U��VW�}�ǃ� ��  H��  H��  H�I  H��  �M�ESj Z�r  �0;1t|�0�+�t3ۅ��Í\�����i  �p�Y+�t3ۅ��Í\�����H  �p�Y+�t3ۅ��Í\�����'  �p�Y+�t3ۅ��Í\����3����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3����r  �p;qt~�p�Y+�t3ۅ��Í\�����I  �p	�Y	+�t3ۅ��Í\�����(  �p
�Y
+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����w  �p�Y+�t3ۅ��Í\����3����R  �p;qt~�Y�p+�t3ۅ��Í\�����)  �p�Y+�t3ۅ��Í\�����  �p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\����3�����  �p;qt~�p�Y+�t3ۅ��Í\������  �p�Y+�t3ۅ��Í\�����x  �p�Y+�t3ۅ��Í\�����W  �p�Y+�t3ۅ��Í\����3����2  �p;qt~�p�Y+�t3ۅ��Í\�����	  �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\������   �p�Y+�t3ۅ��Í\����3�����   �p;qtr�p�Y+�t3ۅ��Í\����u}�p�Y+�t3ۅ��Í\����u`�p�Y+�t3ۅ��Í\����uC�p�Y+�t3ۅ��Í\����3���u"��+�;�������σ���  �$�g����  �P�;Q�tq���Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����u��p��Q�+�t3҅��T����3����v����P�;Q�t}���Q�+�t3҅��T�����N����p��Q�+�t3҅��T�����-����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����}����p��Q�+�t3҅��T����3����X����P�;Q�t}���Q�+�t3҅��T�����0����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T�����^����p��Q�+�t3҅��T����3����9����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�to���Q�+�t3҅��T���u6�p��Q�+�t3҅��T���u�p��Q�+�t3҅��T���t����@��I�+�t3Ʌ����L	����3���u3�[�S  �P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����n����p��Q�+�t3҅��T�����M����p��Q�+�t3҅��T�����,����p��Q�+�t3҅��T����3��������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����x����P�;Q�t}���Q�+�t3҅��T�����P����p��Q�+�t3҅��T�����/����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3����Z����P�;Q�t~�Q��p�+�t3҅��T�����1����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����`����p��Q�+�t3҅��T����3����;����I��@�+�� ���3Ʌ����L	���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����b����p��Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����l����P�;Q�t}���Q�+�t3҅��T�����D����p��Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����s����p��Q�+�t3҅��T����3����N����P�;Q�t~�Q��p�+�t3҅��T�����%����Q��p�+�t3҅��T���������Q��p�+�t3҅��T����������Q��p�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T����3����/���f�P�f;Q�������Q��p�+������3҅��T����  �����P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3����i����P�;Q�t}���Q�+�t3҅��T�����A����p��Q�+�t3҅��T����� ����p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T�����p����p��Q�+�t3҅��T����3����K����P�;Q�t}���Q�+�t3҅��T�����#����p��Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t~�Q��p�+�t3҅��T����������p��Q�+�t3҅��T�����r����p��Q�+�t3҅��T�����Q����p��Q�+�t3҅��T����3����,����P�;Q�t}���Q�+�t3҅��T���������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����������p��Q�+�t3҅��T����3���������P�;Q�t}���Q�+�t3҅��T�����u����p��Q�+�t3҅��T�����T����p��Q�+�t3҅��T�����3����p��Q�+�t3҅��T����3��������p��Q�+������3҅��T���������������M�u��+�t3҅��T�����   �A�V+�t3҅��T�����   �A�V+�t3҅��T�����   �A�N+���   3Ʌ����L	����   �M�u��+�t3҅��T���uh�A�V+�t3҅��T���uK�A�N랋M�u��+�t3҅��T���u �A�N�p����E�M� �	�_���3�_^]���'��kw�
����	
l�LXy	��� ��N�. :[������<��<���������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U�����ISV�uW3��E��}�}��}��FFf�> t����at8��rt+��wt�M��WWWWW�    �������3��S  �  �3ۃM��	�	  �M�3�AFF�f;���  � @  ;��   ����S��   ��   �� ��   ��tVHtG��t1��
t!���u���9}���   �E�   ����   �ˀ   �   ��@��   ��@�   �E�   �   ����   �E����������   �E��}9}�ur�E�   �� �l��TtX��tCHt/��t��������� �  uC��E9}�u:�e������E�   �09}�u%	U��E�   ��� �  u�� �  ��   ��t3���FF�f;������9}���   �FFf�> t�jVh����:  �����`���j ��X�FFf9t�f�>=�G���FFf9t�jh��V�:  ����u��
��   �Djh��V��9  ����u����   �%jh��V��9  �������������   �FFf�> t�f9>�����h�  �u�ES�uP�}8  ����������E�$D�M��H�M�x�8�x�x�H_^[��jhX�Hg��3�3��}�j�C\��Y�]�3��u�;5 [��   � K��9t[� �@��uH� �  uA�F���w�FP�>[��Y����   � K�4�V��i��YY� K���@�tPV�Dj��YYF둋��}��h��j8����Y� K�� K�9tIh�  � �� P��	  YY��� Ku�4�7���Y� K����� P�(�� K�<�}�_;�t�g �  �_�_��_�O��E������   ���nf��Ë}�j�MZ��Y�SVW�T$�D$�L$URPQQh�d�5    �'3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�R  �   �C�d  �d�    ��_^[ËL$�A   �   t3�D$�H3��`���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�  3�3�3�3�3���U��SVWj j hSQ�]  _^[]�U�l$RQ�t$������]� ��U����u�M��*����E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U��3�@�} u3�]�U��SVWUj j h��u�]  ]_^[��]ËL$�A   �   t2�D$�H�3�� ���U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�d�5    �'3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�u�Q�R9Qu�   �SQ� 7�SQ� 7�L$�K�C�kUQPXY]Y[� ����������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �������U��W�}3�������ك��E���8t3�����_�Ë�U���SV�u�M��*����]�   ;�sT�M胹�   ~�E�PjS�����M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�h���YY��t�Ej�E��]��E� Y���E��� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�;
����$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=D? u�E�H���w�� ]�j �u�����YY]Ë�U���(�'3ŉE�SV�uW�u�}�M�������E�P3�SSSSW�E�P�E�P�>?  �E�E�VP�4  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[������Ë�U���(�'3ŉE�SV�uW�u�}�M��0����E�P3�SSSSW�E�P�E�P�>  �E�E�VP�E9  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�0����Ë�U��MSV�u3�W�y;�u��C��j^�0SSSSS�H��������   9]v݋U;ӈ~���3�@9Ew�C��j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W����@PWV������3�_^[]Ë�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���H���u��P������Ɂ���  �P���t�M�_^f�H[�Ë�U���0�'3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��bC  �uЉC�E։�EԉC�E�P�uV������$��t3�PPPPP�V������M�_�s^��3�[�$�����������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j聋��YË�U��E�M%����#�V������t1W�}3�;�tVV�0L  YY��@��j_VVVVV�8��������_��uP�u��t	� L  ����K  YY3�^]Ë�U��E��H]�jhx�\���e� �u�u�$��E��/�E� � �E�3�=  �����Ëe�}�  �uj����e� �E������E��\���������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h�h�wd�    P��SVW�'1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh���Z��3ۉ]�j��O��Y�]�j_�}�;= [}W����� K�9tD� �@�tP�`���Y���t�E��|(� K��� P�$�� K�4�1���Y� K�G��E������	   �E��Z���j�}N��YË�U����UV�uj�X�E�U�;�u� >���  ��=��� 	   ����  S3�;�|;5�Ir'��=����=��SSSSS� 	   �#���������Q  ����W�<� J�����ƊH��u�=����v=��� 	   �j�����wP�]�;��  ����  9]t7�@$����E���HjYtHu���Шt����U�E�E��   ���Шu!�$=����
=���    SSSSS�q������4����M;�r�E�u�R��Y�E�;�u��<���    ��<���    ����h  jSS�u�^  ��D(�E���T,���AHtt�I��
tl9]tg��@�M�E�   �D
8]�tN��L%��
tC9]t>��@�M�}��E�   �D%
u$��L&��
t9]t��@�M�E�   �D&
S�M�Q�uP��4�ؠ���{  �M�;��p  ;M�g  �M��D� ���  �}��  ;�t�M�9
u��� ��]�E�É]�E�;���   �M�<��   <t�CA�M�   �E�H;�s�A�8
u
AA�M�
�u�E�m�Ej �E�Pj�E�P��4�ؠ��u
�L���uE�}� t?��DHt�}�
t����M��L�%;]�u�}�
t�jj�j��u�  ���}�
t�C�E�9E�G������D� @u����C��+E�}��E���   ����   K���xC�   3�@�����;]�rK�@��07 t�����07��u�}:��� *   �zA;�u��@���AHt$C���Q|	���T%C��u	���T&C+���ؙjRP�u��  ���E�+]���P�uS�u�j h��  �l��E���u4�L�P�":��Y�M���E�;EtP�����Y�E�����  �E��  �E��3�;�����E��L0��;�t�M�f�9
u��� ��]�E�É]�E�;���   �E�f����   f��tf�CC@@�E�   �M����;�s�Hf�9
u���Ej
�   �M�   �Ej �E�Pj�E�P��4�ؠ��u
�L���u[�}� tU��DHt(f�}�
t�jXf���M��L��M��L%��D&
�*;]�uf�}�
t�jj�j��u�|  ��f�}�
tjXf�CC�E�9E�������t�@u��f� f�CC+]�]������L�j^;�u�v8��� 	   �~8���0�i�����m�Y����]��\���3�_[^��jh��~T���E���u�F8���  �+8��� 	   ����   3�;�|;�Ir!�8���0�8��� 	   VVVVV�j������ɋ����� J��������L9��t�����;M�Au��7���0�7���    �P��  Y�u���D8t�u�u�u�~������E���7��� 	   �7���0�M���E������	   �E���S����u�  YË�U��QQ�EV�u�E��EWV�E���  ���Y;�u�$7��� 	   �ǋ��J�u�M�Q�u�P�ܠ�E�;�u�L���t	P�7��Y�ϋ����� J�����D0� ��E��U�_^��jh���R������u܉u��E���u�6���  �6��� 	   �Ƌ���   3�;�|;�Ir!�6���8�w6��� 	   WWWWW��������ȋ����� J��������L1��u&�P6���8�66��� 	   WWWWW������������[P�=  Y�}���D0t�u�u�u�u�������E܉U����5��� 	   ��5���8�M���M���E������   �E܋U��?R����u�z  YË�U��E���u�5��� 	   3�]�V3�;�|;�Ir�5��VVVVV� 	   �������3���ȃ����� J���D��@^]Ë�U����'3ŉE�V3�9508tO�=\:�u�C  �\:���u���  �pV�M�Qj�MQP�0���ug�=08u��L���xuω508VVj�E�Pj�EPV�,�P�h��\:���t�V�U�RP�E�PQ�(���t�f�E�M�3�^��������08   ���U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M������E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�l����E�u�M;��   r 8^t���   8]��e����M��ap��Y����3��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�l����:���뺋�U��j �u�u�u�������]Ë�U��EVW��|Y;�IsQ���������<� J����<�u5�=8?S�]u�� tHtHuSj��Sj��Sj��4���3�[���2��� 	   ��2���  ���_^]Ë�U��MS3�;�VW|[;�IsS������<� J�������@t5�8�t0�=8?u+�tItIuSj��Sj��Sj��4����3���e2��� 	   �m2������_^[]Ë�U��E���u�Q2���  �62��� 	   ���]�V3�;�|";�Is�ȃ����� J����@u$�2���0��1��VVVVV� 	   �]���������� ^]�jh�N���}����������4� J�E�   3�9^u6j
��B��Y�]�9^uh�  �FP�#���YY��u�]��F�E������0   9]�t���������� J�D8P�(��E���M���3ۋ}j
�A��YË�U��E�ȃ����� J���DP�,�]�jh8�DM���M��3��}�j�zA��Y��u����b  j�)B��Y�}��}؃�@�<  �4� J����   �u��� J   ;���   �Fu\�~ u9j
��A��Y3�C�]��~ uh�  �FP����YY��u�]���F�e� �(   �}� u�^S�(��FtS�,���@낋}؋u�j
�@��YÃ}� u��F��+4� J��������u�}��uyG�+���j@j ����YY�E���ta�� J���I ���   ;�s�@ ���@
�` ��@�E������}�����σ����� J�DW�����Y��u�M���E������	   �E��L���j��?��Y��������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U��E��H]Ë�U����u�M��%����E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�v  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�O  �EPSj �u�H��M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�}  Y����  �t�Etj�c  Y����v  ����   �E��   j�A  �EY�   #�tT=   t7=   t;�ub��M����@9��{L�H��M�����{,�@9�2��M�����z�@9���M�����z�09��09��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�x  �M��]�� �����������}�E���0��S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj��  Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}�")��� "   ]��)��� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���H8;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P���������uV�,���Y�E�^�Ë�L8�h��  �u(�  �u�����E ���Ë�U��=@8 u(�u�E���\$���\$�E�$�uj�/�����$]���'��h��  �u� !   �J  �EYY]Ë�S��QQ�����U�k�l$���   �'3ŉE��s �CP�s��������u"�e���CP�CP�s�C �sP�E�P�I������s�p������=@8 u+��t'�s �C���\$���\$�C�$�sP�r�����$�P�����$��  �s �  �CYY�M�3��T�����]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj���  f;�u�E�� u9Utj��3�]Ë�U�����U����Dz3��   �U3����  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������"Q���EQQ�$����������  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��#E�����E�m�E��Ë�U��QQ�M��t
�-X9�]���t����-X9�]�������t
�-d9�]����t	�������؛�� t���]����jh`�RA��3�9D[tV�E@tH9p9t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%p9 �e��U�E�������e��U�2A��Ë�U���SVW�����e� �=�H ����   h���8������*  �5|�h��W�օ��  P����$��W��H��P����$��W� I��P�����$��W�I��P����Y�I��thx�W��P����Y�I�I;�tO9ItGP����5I�����YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9� I;�t0P����Y��t%�ЉE���t�I;�tP���Y��t�u��ЉE��5�H���Y��t�u�u�u�u����3�_^[�Ë�U��MV3�;�|��~��u�4?�(�4?�4?��#��VVVVV�    �z��������^]á'��3�9I����Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v�"��j^SSSSS�0�
��������V�u�M��3����E�9X��   f�E��   f;�v6;�t;�vWSV�-������O"��� *   �D"��� 8]�t�M��ap�_^[��;�t2;�w,�$"��j"^SSSSS�0������8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�h�;�t9]�^����M;�t����L���z�D���;��g���;��_���WSV�V������O�����U��j �u�u�u�u�|�����]Ë�U����u�M�������u�u�u�u�<��}� t�M��ap��Ë�U��QQ�'3ŉE��IS�<�VW3�3�G;�u,VVWV�Ӆ�t�=I�/�L���xu
jX�I��I����   ;���   ;�u#9uu�E� �@�EVV�u�u�ӋȉM�;�u3��   ~Ej�3�X���r9�D	=   w�� ����;�t����  ���P�����Y;�t	� ��  �����3�;�t��u�W�u�u�Ӆ�t VV9uuVV��u�uj�WV�u�h���W裻��Y����u�u�u�u���e�_^[�M�3������Ë�U����u�M�臻���u�E��u�u�u�uP�������}� t�M��ap��Ë�S��QQ�����U�k�l$���   �'3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|������������uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�v�����h��  ��x��������>YYt�=@8 uV����Y��u�6�F���Y�M�_3�^襹����]��[Ë�U��UV�uW��H�F��w�� �
�y�B��w�� ��t;�t�_+�^]Ë�U���S�u�M��ѹ��3�9]u.���SSSSS�    �z�����8]�t�E��`p������   W�};�u+����SSSSS�    �D�����8]�t�E��`p������U�E�9XuW�u�:���YY�4V�E� �M�QP�����E����M�QP�������G;�t;�t�+���^8]�t�M��ap�_[�Ë�U��V3�95D?u09uu�D��VVVVV�    �����������9ut�^]����V�u�u�������^]Ë�U���S3�VW9]��   �u�M�蝸��9]u.����SSSSS�    �H�����8]�t�E��`p������   �};�t˾���9uv(���SSSSS�    �	�����8]�t�E��`p����`�E�9Xu�uW�u�A+  ��8]�tD�M��ap��;�E� �M�QP�����E����M�QP������G�Mt;�t;�t�+����3�_^[�Ë�U��V3�95D?u99uu� ��VVVVV�    �g����������'9ut܁}���w�^]�*  V�u�u�u������^]Ë�U��QSV��3�;�u���j^SSSSS�0���������   W9]w���j^SSSSS�0����������   3�9]���A9Mw	�U��j"�ЋM�����"w��]���9]t�-�N�E�   �؋�3��u��	v��W���0�A�E�3�;�v�U9U�rڋE�;Er�럈I���I�G;�r�3�_^[�� ��U��}
�Eu
��}jj
�j �u�u�M�����]Ë�U���4S3��E�VW���]��]��E�   �]�t	�]��E��
�E�   �]��E�P�,  Y��tSSSSS�������M� �  ��u�� @ u9E�t�M������+ú   ��   �tGHt.Ht&�:��������j^SSSSS�0�������  �U����t��   u��E�   @��}��EjY+�t7+�t*+�t+�t��@u�9}����E���E�   ��E�   ��E�   ��]��E�   #¹   ;��   ;t0;�t,;�t=   ��   =   �@����E�   �/�E�   �&�E�   �=   t=   t`;������E�   �E�E�   ��t�(D��#M��x�E�   �@t�M�   �M�   �M��   t	}�� t�M�   ��E�   릨t�M�   ��������u�����������    �   �E�=@�S�u��    �u�E�P�u��u��u�׉E���um�M��   �#�;�u+�Et%�e����S�u�E��u�P�u��u��u�׉E���u4�6������ J�����D0� ��L�P�B��Y���� �u  �u����;�uD�6������ J�����D0� ��L���V����Y�u�� �;�u������    룃�u�M�@�	��u�M��u��6�I�����Ѓ����� JY��Y�M����L��Ѓ����� J���D$� ��M��e�H�M���   �����  �Etrj���W�6�I�����E�;�u�=���8�   tN�6�>M�������j�E�P�6�]����������uf�}�u�E�RP�6�"&  ��;�t�SS�6�%I����;�t��E���0  � @ � @  �}u�E�#�u	M�	E�E#�;�tD=   t)= @ t"=   t)= @ t"=   t= @ u�E���M�  #�;�u	�E���]��E   ��  �E�@�]���  �E��   �#�=   @��   =   �tw;���  �E�;��y  ��v��v0���f  �E�3�H�&  H�R  �E���  �E�   �  jSS�6�������t�SSS�6�n���#���������j�E�P�6����������t�����tk����   �}�﻿ uY�E���   �E�;���   ���b������P���jSS�6���������C���SSS�6�������#����   �����E�%��  =��  u�6�3K��Y�
��j^�0���d  =��  uSj�6�7G�������������E��ASS�6�G������E�﻿ �E�   �E�+�P�D=�P�6�sA������������9}�ۋ������ J�����D$�2M���0������� J�����D$�M�������
ʈ8]�u!�Et��ȃ����� J���D� �}��   ���#�;�u|�Etv�u�� �S�u�E�jP�u������W�u�@����u4�L�P�����ȃ����� J���D� ��6�����Y�����6������ J�������_^[��jh���/��3��u�3��};���;�u�q��j_�8VVVVV�ٺ�������Y��3�9u��;�t�9ut�E%������@tu��u�u�u�u�E�P���i������E��E������   �E�;�t���/���3��}9u�t(9u�t����������� J�D� ��7����YË�U��j�u�u�u�u�u������]Ë�U���SV3�3�W9u��   �];�u"���VVVVV�    �����������   �};�t��u�M������E�9pu?�f��Ar	f��Zw�� ���f��Ar	f��Zw�� CCGG�M��tBf��t=f;�t��6�E�P�P��#  ���E�P�P��#  ��CCGG�M��t
f��tf;�t�����+��}� t�M��ap�_^[�Ë�U��V3�W95D?u3�9u��   �};�u���VVVVV�    ������������`�U;�t��f��Ar	f��Zw�� ���f��Ar	f��Zw�� GGBB�M��t
f;�tf;�t�����+��V�u�u�u�w�����_^]Ë�U��} u3�]ËU�M�Mt�f��tf;uAABB����
+�]Ë�U����  ��f9Eu�e� �e�   f9Es�E��'f�Af#E���E��@�u�M��K����E��p�p�E�Pj�EP�E�jP�#  ����u!E��}� t�E�`p��E��M#��Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���50:N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�,:��+0:;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�50:N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��4:A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;(:�4:��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�(:�<:�3�@�   �<:�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+4:��M���Ɂ�   �ً8:]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5H:N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�D:��+H:;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5H:N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��L:A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;@:�L:��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�@:�T:�3�@�   �T:�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+L:��M���Ɂ�   �ًP:]���@u�M�U�Y��
�� u�M�_[�Ë�U���|�'3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u���SSSSS�    ������3��N  �U�U��< t<	t<
t<uB��0�B���/  �$��[�Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P�x  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �"  =�����.  ��:��`�E�;���  }�ع0<�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��K
3��E��EԉE؉E܋E΋��  3�#�#ʁ� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uB�E����u9u�u9u�u3�f�E���  f;�u!B�C���u9su93u�ủuȉu���  �u��}��E�   �E��M���M���~R�DĉE��C�E��E��M��	� �e� ���O��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?�����  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋M��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9M�w�Mԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�B�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�U�f�EċE؉EƋE܉E�f�U��3�f�����e� H%   � ���e� �Ẽ}� �<����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[�=����Ð�UVnV�V�VW2W�WxW�W�W�W��U���t�'3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�f��t�C-��C �u�}�f��u/��u+��u'3�f;�����$ f��C�C�C0�S3�@�  ��  f;���   3�@f��   �;�u��t��   @uh���Qf��t��   �u��u;h���;�u0��u,h���CjP�&�����3���tVVVVV��������C�*h���CjP�������3���tVVVVV�Σ�����C3��q  �ʋ�i�M  �������Ck�M��������3���f�M��:�ۃ�`�E�f�U�u�}�M�����  }�0<�ۃ�`�E�����  �E�T�˃������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE��P
3ɉM��M��M�M��M��3�� �  �u���  #�#֍4
����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��{����M�����?  ��  f;���  �E�3҉U��U��U�U��U��ɋ�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��V���3�3�f9u���H%   � ���E��\���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �^�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[�%����À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95D[��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E�����Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��3�PPjPjh   @h���D��\:á\:V�5 ����t���tP�֡X:���t���tP��^��U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U���SVW3�jSS�u�]��]��[����E�#��U���tYjSS�u�?�����#ʃ����tA�u�}+����   ;���   �   Sj�L�P�`��E���u�G����    �<���� _^[��h �  �u�  YY�E���|
;�r�����P�u��u��������t6�+��xӅ�wϋu��u��u��   YY�u�j �L�P�P�3��   ������8u�����    ����u��;�q|;�skS�u�u�u�D���#�����D����u�-���YP�H������H��E�#U���u)�[����    �c������L���u�#u��������S�u��u��u�ٷ��#���������3��������U��S�]V�u������ J������0�A$�W�y����   ���� @  tP�� �  tB��   t&��   t��   u=�I��
�L1$��⁀���'�I��
�L1$��₀���a��I��
�L1$�!���_^[u� �  ]����% �   @  ]Ë�U��EV3�;�u�C���VVVVV�    誕����jX�
��I�3�^]Ë�U����  �ȃ�f9M��   S�u�M�諉���M�Q3�;�u�E�H�f��w�� ���aV�   ��f9u^s)�E�Pj�u����������Et9�M싉�   f����q�M�jQj�MQPR�E�P�*  �� ���Et�E�8]�t�M�ap�[�Ë�U����u�M������}�}3���u�u�u�u���}� t�M��ap��Ë�U����'3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[葆���Ë�U����u�M�������E��~�M��Jf�9 t	AA��u���+�H�u �uP�u�u�u�p��}� t�M��ap����%0������̋M��8����M����]����T$�B�J�3��������饂���M��
����M����/����T$�B�J�3��څ�����w����M��\P���M��ԟ���M��̟���M��DP���M��<P���M�鴟���M�鬟���M�餟��h�h�   h�=�E�P�L�����ËT$�B�J�3��c����@�� ����M���O����l�����O���M���O���M��ڰ���M��B����M��O���M��2����M��O����l����O����4����O����P����O���M��O���M�������M������M������M������M��ٞ���M��QO���M��ɞ���M�������M�鹞���M�鱞���M�驞���M�類���T$�B��0���3��y�����������M������M��s����M���N���T$�B�J�3��F�����������M��H���h�h�   h�=�EP��������h�h�   h�=��H���P�р����ÍM������M�������E����   �e���M�����ÍM��ܝ���M��ԝ���T$�B��D���3�謃������I��������̍M��(����M��п���T$�B�J�3��{����h������M�������M�饿���E����   �e���M�]���ËT$�B�J�3��7�����������M�鹯���M��a����T$�B�J�3������������M�鎯���E����   �e���M��&���ËT$�B�J�3��Ђ�����m���M��R����M�������T$�B�J�3�襂���@��B���M��'����M��Ͼ���E����   �e���M�M��ËT$�B�J�3��a����|���~���M�c����T$�B�J�3��>��������~���M��@����T$�B�J�3���������~���E����   �e���M����ÍM������M�������M��������p��������M�������P����֛���M��Λ���M��ƛ���M�龛����`���鳛����@���騛���M�頛���T$�B��@���3��x�������~���M��*����M��������M���0�����M���H�	����M���`������M���x�����M����   �����M����   �׬���T$�B�J�3���������}���M�鴬���M���马���M���0鞬���M���H铬���M���`鈬���M���x�}����M����   �o����M����   �a����T$�B�J�3�茀������)}���M�鎚����|���郚��������x�����<����m����M��e����M��]����M��U�����\����J����M��B����M��:�����L����/�����l����$�����,����������������������������������������������������������M��ڙ���M��ҙ����l����Ǚ����L���鼙���M�鴙���T$�B������3�����L��)|��������鋙�������這���������u�����(����j����M��b����������W�����x����L����������A����������6�����(����+��������� ���������������x����
�����H����������H����������h���������X����ޘ����x����Ә���������Ș���M������������鵘����X���骘����h���韘��������锘��������鉘���������~����������s���������h����������]����������R����������G�����h����<����M��4����M��,���������!�����x������������������������ ������������������������������ߗ����8����ԗ����X����ɗ����h���龗���M�鶗���M�鮗����(���飗����H���阗����8���鍗��������邗���������w����������l����������a����������V���������K�����8����@�����X����5����M��-����M��%�������������������������8��������T$�B��T���3���|���H��yy���M��ޖ����\����SG����0����HG���M�������M�鸖���M�鰖����0����%G���M�靖���M�镖���M�鍖���M�酖���M��}����M��u����M��m����M��e����M��]����M��U����M��M����M��E�����L����:�����x����/����M��'����M������� ��������� ����	��������������M��������<��������M�������h����ؕ���M��Е���M��ȕ���M�������� ���鵕����<���骕����h���韕���T$�B������3��w{���|��x���M�y�����`����n����M��f����M��^����M��V�����p����K����M��C����M��;�����P����0�����4����%��������������������������������������������(����nE����D����cE���M��[E���M��SE���M��˔���M��Ô���M�黔���M�鳔���M�體���M�飔���M�雔���T$�B������3��sz������w���M���D���M��m����M��e�����D�����D����D�����D���M��G����M��?����M������M��/�����p����$����M�������P���������4��������M��������`��������M������M������T$�B��0���3��y������Xv���������:D���M�鲓���M�骓����(����D����(����D����`���鉓����������C���M��v����M��n�����(�����C����(�����C����������C���M��E����M��=�����(����C����(����C���M������M������M������M��g���M�����M�������M������M������M��ߒ���M��ג���M��ϒ���M��ǒ���M�鿒���M�鷒�������鬒����`���顒�������閒���M������D���郒���M��{����M��s����M��k���������`�����`����U���������J����M��B����M��:���������/�����`����$�������������������������������������鸴����������������������M��ڑ���M��ґ���������������`���鼑���M�鴑��������驑��������鞑���M�閑���M�鎑��������郑���������x���������m����T$�B��D���3��Ew���`���s����������������̍M��8����E����   �e���M� ���ËT$�B�J�3���v������s�����̋E����   �e���M����ËT$�B�J�3���v������_s�������������̍M鸐���M�������T$�B�J�3��v������(s���M������M��A���T$�B�J�3��`v��� ���r���M��b����M��ڢ���M�邲���M��ʢ���M��¢���M��j����M��b����M��@���T$�B�J�3��v���D��r���M������M������M��'����M��o����M��g����M������M������M��O@���T$�B�J�3��u������Gr���M�鬏���M��$����M��̱���M������M������M�鴱���M������M�������M�霱���M���?���T$�B�J�3��?u������q���M��A����M�鹡���M��a����M�驡���M�顡���M��I����M��A����M�鉡���M��1����M��y?���T$�B�J�3���t������qq����4����ӎ����4����Ȏ�������齎�������鲎�������駎����$���霎����@���鑎���� ���醎����0����{���������������T$�B�����3��Ht���J�3��>t�������p���M��@����T$�B�J�3��t���p��p���M��m���M���$�>���M���@�>���M���\�|>���M����   龘���T$�B�J�3���s������fp���M�����M��$�@>���M��@�5>���M��\�*>���M���   �l����M���   �>����T$�B�J�3��is������p����0����8����������]����������R����������G���������<����� ����1����������&����T$�B������3���r���J�3���r���4��o���������õ��������������p����݌����`����Ҍ����(����ǌ���� ���鼌�������鱌����`���馌����p���雌�������鐌���� ���酌����(����z�����p����o����������d����������Y�����D���������4����C�����`����8�����p����-���������"����� ���������(���������`���������p������������������� ����������(����Ջ����p����ʋ����`���鿋����8���鴋��������驋��������鞋����8���铋��������鈋���������}����T$�B������3��Uq���J�3��Kq�������m���E���   �e���M�}���ÍM��Ă���M�鼂���T$�B�J�3��q������m���������F����������;����������������d���������T����ڊ���������ϊ����(����Ċ����D���鹊����d���鮊����T���飊��������阊����(���鍊����D���邊����l����w����������l�����t�����:����t�����:���������K�����t����Ё����l���饁���������Z�����D���������P���餁����l����y����������.�����x����3����T$�B��L���3���o���J�3���o�����^l�������������������鵉��������骉��������韉���������:���������	:���������~����������s�����������9����������9���������"����������G����������<����������1����������&���������������d������������������������������d������������������������و���������Έ����t����È��������鸈����T���魈����D���颈���T$�B������3��zn���J�3��pn�����k�����������̋M��h����M���L�]����M���\�R����M���p�G����T$�B�J�3��"n���(��j�������������̋M������M���L�����M���\�����M���p������T$�B�J�3���m���l��oj�������������̋M���e���T$�B�J�3��m������=j�����������̋M���H��^���T$�B�J�3��pm�����j�����������̋T$�B�J�3��Km���|���i������̋EP�M�Q�S�����ËT$�B�J�3��m�����i�����̋M���i���T$�B�J�3���l���0��i��������������̋EP�M�Q������ËT$�B�J�3��l������Wi�����̋M��8`���M����=~���M��� �2~���M���<�'~���M���X�~���T$�B�J�3��gl������i��̋M���_���M�����}���M��� ��}���M���<��}���M���X��}���T$�B�J�3��l��� ��h��̍M��}���T$�B�J�3���k���J�3���k���T��h����̍M��x}���T$�B�J�3���k���J�3��k������Vh����̋M��nt���T$�B�J�3��k������0h��������������̋EP�e��YËE����   �e���M���|��ËT$�B��\���3��Dk�������g���������������̍M���|���T$�B�J�3��k���J�3��	k�����g����̍M��|���T$�B�J�3���j������g��������������̍M��X^���T$�B�J�3��j������Pg��������������̋E�P�d��YËE����   �e���M��|��ËT$�B��\���3��dj���8��g���������������̋EP�M�Q�c�����ËT$�B�J�3��*j�������f�����̍M��{���M��{����l����{���T$�B��t���3���i������f��������̋M��r���T$�B�J�3���i���X �`f��������������̋M��f���T$�B�J�3��i���� �0f��������������̍M��x���T$�B�J�3��ci���� � f��������������̋T$�B��l���3��8i���J�3��.i�����e���������̍�L����E\���������:\���T$�B������3���h�����e�������������̋EP�M�Q������ËT$�B�J�3��h���8�We�����̋M��s���T$�B�J�3��h���d�0e��������������̋M���P��Y���T$�B�J�3��`h������d�����������̍M�x[���T$�B�J�3��3h������d��������������̍M����T$�B�J�3��h�����d��������������̍M��y���E�P�M�Q�������ËT$�B�J�3���g���J�3��g���P�Ud���̍M����T$�B�J�3��g�����0d��������������̋M��8d���T$�B�J�3��cg����� d��������������̋E����   �e���M��X�uX��ËM���yX���T$�B�J�3��g���0�c���������������̋E����   �e���M��P�%X��ËM���)X���T$�B�J�3���f���l�ac���������������̍M��hc���T$�B�J�3��f�����0c��������������̍M��8c���M��p ���T$�B�J�3��[f���,��b������̍M���w���M���w���T$�B�J�3��+f���J�3��!f�����b������������̋M����w���T$�B�J�3���e���,�b�����������̍M,�|���M�|���T$�B�J�3��e���`�Xb������̍M,��{���M��{���M���{���T$�B�J�3��e����� b��������������̋M��ؼ���T$�B�J�3��Se������a���������������hȪjh�=�E�P��a����ËM��/���T$�B�J�3��
e�����a���M��X���T$�B�J�3���d���(�a���M�������T$�B�J�3���d���T�aa���M������M����Kv���T$�B�J�3��d�����3a���M��X���u��^��YËT$�B�J�3��id�����a���M���u���T$�B�J�3��Fd������`���T$�B�J�3��+d����
��`�������h`�輈��Yù`>�W��h��覈��Y�h��蚈��Yù?��V��hɒ脈��Y�hӒ�x���YÃ=�= uK��=��t��=�Q<P�B�Ѓ���=    ��=��tV��� .��V�]������=    ^ù`>�V����>�g����?�V���?�^��                                                                                                                                                                                                                                                                                                   4 B R b t � � � �  ( @ X d x � � � � � �   , > J Z p � � � � � � � � � 
    2 F T b p � � � � � � � � �   0 > T n � � � � � �    2 D V l � � � � � �    " 0 > N     �         �>�T��2�        i}Z]2y��        �i�y                    �4LM          �� �� bad allocation  x� " � p ��@  �� ` �[3D-COAT     c:\program files\maxon\cinema 4d r11.5\plugins\applink_3dcoat\source\applinkdialog.cpp  Start import!   To import a new object? File exists!    export.txt  Folder ..\MyDocuments\3D-CoatV3\Exchange not found! 3D-CoatV3   Exchange    preference.ini  3D-Coat.exe is run! 3D-Coat.exe not found!  open        c:\program files\maxon\cinema 4d r11.5\plugins\applink_3dcoat\source\applinkexporter.cpp    
   c:\program files\maxon\cinema 4d r11.5\resource\_api\ge_dynamicarray.h  ]   autopo  curv    prim    alpha   vox retopo  ref uv  ptex    mv  ppp [   # end   v       # begin      vertices
            �?vt   texture vertices
  /   f   usemtl   faces
 g   mtllib  mtl map_    illum 2
    Tr 0.000000
    Ns 50.000000
   Ks  Kd  Ka 0.300000 0.300000 0.300000
  newmtl  No selected objects!    Object "    " has no UVW tag.
UV coordinates can't be exported. Material not found on   object. Default Name    Export object   #Cinema4D Version:  %d.%m.%Y  %H:%M:%S  #File created:  #Wavefront OBJ Export for 3D-Coat
  File     write success!   ��import.txt  output.obj  obj �� � �x��� 0�� ��0� ��� ����  �  � p� P� �� �� �� 0�  � `�           Y@�p� @� @� �� P� �� `� �� `�  �  � �� �� �� \��� �� @� �� �� �� `� �� `�  � P� �� �� �� ���� �� �� �� p� p� �� �� Selection   Error on inserting phongTag. Object:    Create objects...   Memory allocation error for material.   �� P��)P��� ��`� �� `� ��@Pp4��`
�
���
�
4�`
�
���
�
vector<T> too long  bad cast    ios_base::eofbit set    ios_base::failbit set   ios_base::badbit set    ���9    X       P   f   vt  Gathering of data...     not found!  can not removed!   normalmap   displacement %f displacement    map_Ks %s   map_Ks  map_Kd %s   map_Kd  Ke %lf %lf %lf  Ke  Ks %lf %lf %lf  Ks  Ka %lf %lf %lf  Ka  Kd %lf %lf %lf  Kd  illum %d    illum   d %lf   d   Ns %lf  Ns  newmtl %s    open!      c:\program files\maxon\cinema 4d r11.5\plugins\applink_3dcoat\source\applinkimporter.cpp    vt %lf %lf %lf  vt %lf %lf  v %lf %lf %lf   g %s    mtllib %s   Parse file...   Open file:  .   textures.txt    ��pN�Lp� ���0�P�@�icon_coat.tif   c:\program files\maxon\cinema 4d r11.5\plugins\applink_3dcoat\source\applinkpreferences.cpp          �f@-DT�!	@      �?������������ ��Ѕ�[     @�@������������ ��Ѕ �H�p�����0�@��� �P� �`�0�c:\program files\maxon\cinema 4d r11.5\resource\_api\c4d_gui.cpp    ������������ ��Ѕ�    ������������ ��Ѕ0���������Т����@�P� �0�Progress Thread 99% 0%  ~   %   c:\program files\maxon\cinema 4d r11.5\resource\_api\c4d_file.cpp   %s         c:\program files\maxon\cinema 4d r11.5\resource\_api\c4d_string.cpp  B   KB  MB       P? GB     ����MbP?`�`|Pb��@|    c:\program files\maxon\cinema 4d r11.5\resource\_api\c4d_baseobject.cpp ��������p~@����~P� �`�0�      �c:\program files\maxon\cinema 4d r11.5\resource\_api\c4d_resource.cpp   #   M_EDITOR    @���res    ? �Ngm��C   ����AT���� ��    c:\program files\maxon\cinema 4d r11.5\resource\_api\c4d_pmain.cpp  �������^    c:\program files\maxon\cinema 4d r11.5\resource\_api\c4d_libs\lib_ngon.cpp              c:\program files\maxon\cinema 4d r11.5\resource\_api\c4d_basebitmap.cpp �� �c:\program files\maxon\cinema 4d r11.5\resource\_api\c4d_gv\ge_mtools.cpp   ��p�,� �x�����%�*   C   �����g��
string too long invalid string position r            
   !   "   2   *            #   3   +       w   a   r b     w b     a b     r +     w +     a +     r + b   w + b   a + b   \�K���J�J���_��Unknown exception   �����csm�               �                          �?      �?3      3            �      0C       �       ��                                                                                                                                                                                                                                                                                                        ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������LC_TIME LC_NUMERIC  LC_MONETARY LC_CTYPE    LC_COLLATE  LC_ALL  ȹ    ~-��8-~-��8-"��8-y���8-!���8-c�	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ _., _   ;   =   =;  @�'>�bad exception   EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    `?�?e+000          �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    CorExitProcess  m s c o r e e . d l l     �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:    ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx              �������             ��      �@      �              �?5�h!���>@�������             ��      �@      �        HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun united-states   united-kingdom  trinidad & tobago   south-korea south-africa    south korea south africa    slovak  puerto-rico pr-china    pr china    nz  new-zealand hong-kong   holland great britain   england czech   china   britain america usa us  uk  swiss   swedish-finland spanish-venezuela   spanish-uruguay spanish-puerto rico spanish-peru    spanish-paraguay    spanish-panama  spanish-nicaragua   spanish-modern  spanish-mexican spanish-honduras    spanish-guatemala   spanish-el salvador spanish-ecuador spanish-dominican republic  spanish-costa rica  spanish-colombia    spanish-chile   spanish-bolivia spanish-argentina   portuguese-brazilian    norwegian-nynorsk   norwegian-bokmal    norwegian   italian-swiss   irish-english   german-swiss    german-luxembourg   german-lichtenstein german-austrian french-swiss    french-luxembourg   french-canadian french-belgian  english-usa english-us  english-uk  english-trinidad y tobago   english-south africa    english-nz  english-jamaica english-ire english-caribbean   english-can english-belize  english-aus english-american    dutch-belgian   chinese-traditional chinese-singapore   chinese-simplified  chinese-hongkong    chinese chi chh canadian    belgian australian  american-english    american english    american    ��ENU ��ENU ��ENU ��ENA ��NLB t�ENC p�ZHH l�ZHI d�CHS P�ZHH <�CHS (�ZHI �CHT �NLB ��ENU ��ENA ��ENL ��ENC ��ENB ��ENI ��ENJ ��ENZ t�ENS X�ENT L�ENG @�ENU 4�ENU $�FRB �FRC  �FRL ��FRS ��DEA ��DEC ��DEL ��DES ��ENI ��ITS |�NOR h�NOR T�NON <�PTB (�ESS �ESB �ESL ��ESO ��ESC ��ESD ��ESF ��ESE ��ESG x�ESH h�ESM X�ESN D�ESI 4�ESA  �ESZ �ESR ��ESU ��ESY ��ESV ��SVF ��DES ��ENG ��ENU ��ENU ��USA ��GBR ��CHN ��CZE ��GBR |�GBR t�NLD h�HKG \�NZL X�NZL L�CHN @�CHN 4�PRI ,�SVK �ZAF �KOR  �ZAF ��KOR ��TTO ��GBR ��GBR ��USA ��USA 6-0   OCP ACP Norwegian-Nynorsk   c c s   U T F - 8   U T F - 1 6 L E     U N I C O D E    Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   ->* &   +   -   --  ++  ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        p�h�\�P�D�8�,�$�����`�D�0���������������������������������������������������������������������������|�x�t�p�l�`�T�L�@�(�����������h�D�(��������������t�P�H�<�,��������x�L�0��������t���_nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh    GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp       SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    1#QNAN  1#INF   1#IND   1#SNAN  CONOUT$     H                                                           'P�^   RSDS���2��[A��ƬH+��   C:\Program Files\MAXON\CINEMA 4D R11.5\plugins\AppLink_3DCoat\obj\Applink_3DCoatR115_Win32_Release.pdb               ��           ������            ����    @   ��          ����    @   ��           ����                @ �           �(�D�    @        ����    @   �\         ����    @   `�           p�D�                x ��           ����    x         ����    @   ��           ������    �        ����    @   ��           ����    �        ����    @   ��            � D�           T�`�|�    �        ����    @   D��        ����    @   ��           ����    �         ����    @   ��           !��           ��� �x���    !       ����    @   ��L!              P   <�           L�\�`�|�    L!       ����    @   <��               @   D��               @   ��            L!<�            �!��           �������    �!       ����    @   ��            �!(�           8�@�    �!        ����    @   (�            �!p�           ����@�    �!       ����    @   p�            0"��           ��������    0"       ����    @   ��    P       P"�           �4�� �x���    P"       ����    @   �            �"d�           t���@�    �"       ����    @   d�            �"��           ����D�    �"       ����    @   ��             #��           ��D�     #       ����    @   ��             #H�           X�h���D�     #       ����    @   H�            @#��           �����D�    @#       ����    @   ��    X       �#��           ���� �x���    �#       ����    @   ��           <�H�d�    �#       ����    @   ,��#        ����    @   ��           ��d�                �#��           ����H�d�    �#       ����    @   ��              ��            ($�            �,���    ($       ����    @   �            D$\�           l�t�    D$        ����    @   \�            `$��           ������    `$       ����    @   ��            x$��            ������    x$       ����    @   ��           <�D�    �$        ����    @   ,�            �$t�           ����    �$        ����    @   t�            �$��           ����D�    �$       ����    @   ��            %�           �$�t�    %       ����    @   �            �#��            X%h�           x���    X%        ����    @   h�            �%��           ����    �%        ����    @   ��            �%��           ��    �%        ����    @   ��            �%@�           P�\�D�    �%       ����    @   @�            �%��           ����    �%        ����    @   ��            &��           ������    &       ����    @   ��            D& �           0�@���D�    D&       ����    @    �            'p�           ����    '        ����    @   p�            \ `�            d#��           ����D�    d#       ����    @   ��            �'�           (�4�D�    �'       ����    @   �	� � �w � � p Ap �p �q �q lr �r �r s Ks vs �s �s  t �t u �u �v <y �z �{ ]| �~ ! Y � � � q� ܀ G� Ё  � R� �� � Ä � M� �� �� I� {� �� Ј � (� a� �� � (� X� �� Ԋ � 8� h� �� � +� X� �� �� �� &� a� �� �� � � Y� �� �� � W� �� �� �� +� `� �� Ȑ � 4� W� �� �� Ց �                 ���� p    p"�   ��                       ����.p    6p"�   �                       "�	   d�                       ����\p    dp   lp   tp    |p    �p    �p    �p    �p"�   ��                       �����p    �p   �p�����p   �p   �p   q   q   q   !q	   ,q
   7q	   7q   7q   7q   7q   ?q   Gq   Oq   Wq   _q   gq   oq   wq   q   �q   �q   �q�����q    �q   �q"�   ��                       "�	   �                       ����r����3r   ;r����;r   Cr   \r   dr�����q�����q�����r    �r"�   X�                       �����r    �r   �r"�   ��                       �����r    s"�   ��                       ����*s    2s"�   ��                       ����fs    ns"�   0�                       �����s    �s   �s"�   d�                       �����s"�   ��                       �����s"�   ��                       "�   �                       ����t    4t    <t    Dt    Lt    Wt    _t    jt    rt    zt    �t    �t    �t"�   ��                       �����t    �t   �t   �t   �t   �t   �t   u"�   �                       ����4u    <u   Gu   Ru   ]u   hu   su   �u"�   p�                       �����u    �u   �u   �u   �u   �u   �u    �u�����u   �u	   �u
   �u   �u   �u   v   v   v   'v   2v   =v   Hv   Sv   ^v   fv   nv   yv   �v"�B   l�                       �����v    �v   �v   �v   �v   �v   �v    �v�����v   �v	   �v
   �v   �v   
w   w    w   +w   6w   Aw   Lw   Ww   bw   mw   xw   �w   �w   �w   �w   �w   �w   �w   �w   �w    �w!   �w   �w#   x$   x%   x&   x'   *x(   5x)   @x*   Kx+   Vx,   ax-   lx.   wx   �x0   �x1   �x2   �x3   �x4   �x5   �x6   �x7   �x8   �x9   �x:   �x;    y   y=   y>   y?   &y@   1y"�$   ��                       ����Zy    by   my   xy   �y   �y   �y   �y   �y   �y    �y
   �y   �y   �y    �y   �y   �y   �y   �y    �y   z   z   z   !z   ,z   7z   Bz   Jz   Uz   ]z   hz   pz   xz    �z!   �z"   �z"�   ��                       �����z    �z   �z    �z   �z   �z   �z   �z   �z   {	   {
   {   &{   1{   <{   G{   R{   ]{   e{   m{   u{   }{   �{   �{   �{   �{"�   ��                       �����{    �{   �{   �{    �{    �{    �{    |   	|   |	   |
   $|   /|   :|   B|   M|   U|"�?   ��                       ����{|    �|   �|   �|    �|    �|    �|   �|   �|   �|   �|   �|   �|   �|   }   }   }   !}   )}   1}   9}   A}   I}   Q}   Y}   a}   i}   q}   y}   �}   �}   �}   �}   �}!   �}"   �}"   �}$   �}%   �}&   �}'   �}"   �})   �}*   ~+   ~,   ~"   '~.   2~"   =~0   H~1   S~0   y~3   �~4   �~5   �~0   ^~0   f~0   n~0   �~:   �~;   �~<   �~   �~����     "�   |�                       ����@"�   ��                       �����    �"�   ��                       �����    �"�   �                       "�   h�                       ����������   �   �   �   �   �   �"�   ��                       ����1�����9�   A�   I�   Q�   Y�   a�   i�"�
   0�                       ������������   ��   ��   ��   ��   ��   Ā   ̀   Ԁ"�
   ��                       ������������   �   �   �   �   '�   /�   7�   ?�"�
   �                       ����b�����m�����x�������   ��������   ��   ��   ������Ł������"�   h�                       "�   ��                       �����    #�   .�   9�   D�"�   �                       ����m�    u�   ��   ��   ��   ��"�   X�                       ����͂    ؂   �   �   ��   �    �"�#   ��                       ����B�    M�   X�   c�   n�   y�   ��   ��   ��   ��	   ��
   ��   ƃ   у   ܃   �   �   ��   �   �   �   )�   4�   ?�   J�   U�   `�   k�   v�   ��   ��   ��   ��    ��!   �������    �    �"�   ��                       "�   ,�                       ����/�    :�   E�   P�   [�   f�   q�   |�   ��   ��	   ��
   ��   ��   ��   Ʌ   ԅ   ߅   �   ��    �    �   �   �   !�   ,�   ,�   7�   B�"�   0�                       ����u�    ��������   ��   ��������������      ͆����؆�����
   �
   ��   �   �   �   %�
   0�   ;�   F�   Q�   \�
   g�   r�   }�   ��   ������Ї    ؇   �   �"�   �                       ���� �    (�   3�   >�"�   L�                           ��     ��   ����    @     ����        �     \     ����       ������p�"�   ��                       ������"�   �                       @           J@           �����    ����                  "�   \�   ��                           L�              <�@           o             ������        ������    "�   ��   ��               ���� �"�   (�                       @           
             T�����        P�����    "�   x�   d�               "�   ��                       ������    ��   ��   ��   ��"�   $�                       ����Љ    ؉   �   �   ������ �"�   L�                       ����P�"�   x�                       ������"�   ��                       ������    ��������"�   ��                       ���� �"�   �                           �    H�   X�t���     #    ����    (   �"    �"    ����    (   �!����0�"�   ��                           T�    ������`�"�   ��                          ���    d#    ����       7�������    ��������"�    �                       @           y&             \�����        ������    "�   ��   l�                   P     �������������� �"�   ��                           4 ��    @#    ����    (   @(     #    ����    (   �'����P�"�   P                        ������"�   |                        ������"�   �                        @           �,@           �,����    ����    ����    ����    "�   �    8                             �             � @           �0@           z/"�   �   �                             p            `����    ����    �����              �����@           i3             �����        P�����    "�                      ������"�   \                       ������"�   �                       ������"�   �                       �����"�   �                       @           �8            ����@�           H�        "�   0                  @           L;            t"�   �   �               ����������    ����                         ������"�   �                       ������            ��"�                          ����0�            L�"�   T                       @           �@            �"�   �   �               ������                                     @           �B            "�   P                  ������    ��                                     @           �G@           �F"�   �   �                             �            �����    ����    ������              ��������� �"�   $                       ����P�    X�"�   P                       ������    ��   ��"�   �                       ������"�   �                       ���������	�"�   �                       ����,�"�                           ����O�"�   L                       ����r�    z�"�   x                       ������    ��"�   �                       ����͑"�   �                           \�       ,t���    D&    ����    (   ������    ����    ����    I    ����    ����    ����    z    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    u        A����    ����    ����    �    ����    ����    ����    �	    ����    ����    ����    �    ����    ����    ����    /    ����    ����    ����    f    ����    ����    ����    ����    ����    ����    �    ����    ����    ����    �    ����    ����    ����    -    ����    ����    ����    �9        H9        Y9    ����    ����    ����    N:    ����    ����    ����    �?    x?�?����    ����    ����_@h@@           FA����    ����                  �
"�   �
   �
                   ����    ����    ����    ~B    �A�A����    ����    ����eDiD    ����    ����    �����DE    >    |   ���    �'    ����       �I    ����    ����    ����    �L����    �L����    ����    ����    �N����    �N����    ����    �����P�P    ����    ����    ����2Q6Q    ����    ����    ����    S    ����    ����    ����    vV    ����    ����    ����    DZ    ����    ����    ����\�\    ����    ����    ����    8l    ����    ����    ����I~M~    ����    ����    ����    ��    ����    ����    ����    s�    ����    ����    ����    :�    ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    |�    ����    ����    ����    �    ����    ����    ����    X�    ����    ����    ����    ��    ����    ����    ����    I�    ����    ����    ����    q�    ����    ����    ����        ����    ����    ������    ����    ����    ����/    ����    ����    ����    �    ����    ����    ����    �#    ����    ����    ����    ?%    ����    ����    ����    �)    ����    ����    ����    y+        �*����    ����    ����6#6    ����    ����    ����    �G�         �  � ,         � T�                     4 B R b t � � � �  ( @ X d x � � � � � �   , > J Z p � � � � � � � � � 
    2 F T b p � � � � � � � � �   0 > T n � � � � � �    2 D V l � � � � � �    " 0 > N     �     C CloseHandle EProcess32Next Module32First CProcess32First  � CreateToolhelp32Snapshot  KERNEL32.dll  ShellExecuteExA SHELL32.dll �InterlockedIncrement  �InterlockedDecrement  !Sleep �InitializeCriticalSection � DeleteCriticalSection � EnterCriticalSection  �LeaveCriticalSection  �RtlUnwind -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent ZRaiseException  �GetLastError  �HeapFree  � DeleteFileA �GetCurrentThreadId  oGetCommandLineA �HeapAlloc �LCMapStringA  zWideCharToMultiByte MultiByteToWideChar �LCMapStringW  [GetCPInfo �GetModuleHandleW   GetProcAddress  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �SetLastError  RGetACP  GetOEMCP  �IsValidCodePage �GetModuleHandleA  �HeapCreate  �HeapDestroy WVirtualFree TVirtualAlloc  �HeapReAlloc �SetHandleCount  ;GetStdHandle  �GetFileType 9GetStartupInfoA �WriteFile �GetConsoleCP  �GetConsoleMode  AFlushFileBuffers  hReadFile  �SetFilePointer  ExitProcess �GetModuleFileNameA  JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW �GetEnvironmentStringsW  TQueryPerformanceCounter fGetTickCount  �GetCurrentProcessId OGetSystemTimeAsFileTime �HeapSize  �GetLocaleInfoA  =GetStringTypeA  @GetStringTypeW  mGetUserDefaultLCID  � EnumSystemLocalesA  �IsValidLocale �InitializeCriticalSectionAndSpinCount �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW �SetStdHandle  �LoadLibraryA  �GetLocaleInfoW   CreateFileW x CreateFileA �SetEndOfFile  #GetProcessHeap      �4LM    �          � � � P� �   Applink_3DCoatR115.cdl c4d_main                                                                               ̡Ȱ    .?AVApplinkDialog@@ Ȱ    .?AVGeDialog@@  ̡̡Ȱ    .?AVbad_alloc@std@@ Ȱ    .?AVexception@std@@ Ȱ    .?AVfacet@locale@std@@  Ȱ    .?AVcodecvt_base@std@@  Ȱ    .?AUctype_base@std@@    Ȱ    .?AVios_base@std@@  Ȱ    .?AV?$_Iosb@H@std@@ Ȱ    .?AV?$basic_istream@DU?$char_traits@D@std@@@std@@   Ȱ    .?AV?$basic_ios@DU?$char_traits@D@std@@@std@@   Ȱ    .?AV?$ctype@D@std@@ Ȱ    .?AV?$basic_streambuf@DU?$char_traits@D@std@@@std@@     Ȱ    .?AV?$basic_stringbuf@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    Ȱ    .?AV?$codecvt@DDH@std@@ Ȱ    .?AV?$basic_istringstream@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@    Ȱ    .?AV?$basic_filebuf@DU?$char_traits@D@std@@@std@@   Ȱ    .?AVlogic_error@std@@   Ȱ    .?AVruntime_error@std@@ Ȱ    .?AVlength_error@std@@  Ȱ    .?AVfailure@ios_base@std@@  Ȱ    .?AVbad_cast@std@@  Ȱ    .?AV?$basic_ifstream@DU?$char_traits@D@std@@@std@@  ̡̡Ȱ    .?AVCommandData@@   Ȱ    .?AVBaseData@@  Ȱ    .?AVApplinkPreferences@@    ̡̡̡Ȱ    .?AVGeModalDialog@@ Ȱ    .?AVGeUserArea@@    Ȱ    .?AVSubDialog@@ Ȱ    .?AViCustomGui@@    ̡̡̡̡̡̡̡̡̡̡Ȱ    .?AVGeSortAndSearch@@   Ȱ    .?AVNeighbor@@  Ȱ    .?AVDisjointNgonMesh@@  ̡Ȱ    .?AVTexturePreview@@    ̡̡̡̡̡̡̡̡Ȱ    .?AVC4DThread@@ ̡̡̡̡̡̡̡Ȱ    .?AVGeToolNode2D@@  Ȱ    .?AVGeToolDynArray@@    Ȱ    .?AVGeToolDynArraySort@@    Ȱ    .?AVGeToolList2D@@  ̡����̡Ȱ    .?AV_Locimp@locale@std@@    ̡   ̡Ȱ    .?AVout_of_range@std@@  ̡4�t�t�x�|�������������������        ̡
   Copyright (c) 1992-2004 by P.J. Plauger, licensed by Dinkumware, Ltd. ALL RIGHTS RESERVED.      N�@���D̡Ȱ    .?AVtype_info@@             u�  s�          ̡            fmod         ��/�������/���-�-�W�-�����/���sqrt    ����   ��        ̡Ȱ    .?AVbad_exception@std@@ ��������    ̡                                                                                                                                                                                                                                                                                                                                                abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     (�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    ����    C                                                                                              8-            8-            8-            8-            8-                              �6        ����� 6@-   @-(                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                                   K     K                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �����
                                                          �      x   
   ?     �   ��	   ��
    �   ��   ��   ��   t�   <�   �   ܿ   ��   |�   \�   ��    ��!   Ƚ"   (�x   �y   �z   ���   ��   �����               ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      ������������� ����.�3�I�N�j�z���������������.�B�b�g���������������%�*�J�^�v���������������.�N�S�m�r���������������6�J�b�  ����������������������t�l�`�\�X�T�P�L�H�D�@�<�8�4�0�(����L������������������������	          6.   �6�H�H�H�H�H�H�H�H�H�6   .       �                                                                                                                                                                                                                                   �&         ؼ   ܼ   ̼   м   p�   h�!   `�   ļ   ��   ��   X�   P�   ��   ��    ��   ��   ��   H�   ��   @�   8�   0�   (�    �"   �#   �$   �%   �&    �      �      ���������              �       �D        � 0         �p     ����    PST                                                             PDT                                                             �9�9����        ����           ���5      @   �  �   ����             ������������   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
                                                                                                                       �   00A0V0d0�0�0�0�0:1$2M2�2�2�2@3V3m3�3�3�3�344&4>4f4�4�4�4v6�6�6x7�7�7�78�8�8�89|9�9:s:�:�:�:*;@;�<�<�<f=w=�=F>[>�>�>�>�>�>�>|?�?�?�?      �   0)0a0�0�0�0�0	1+151O1f1�1�1d2�2�2�2�4�4535F5^5�5�5�5L6a6u6�6�6�6�6�677r7�7�7�78_8�8�8�89'9~9�9::z:�:�:;;';@;P;_;�;�;�;�;<<'<?<M<\<�<6=J=`=t=�=�=�=�=�=>->G>m>�>�>�>�>?/?W?w?�?�?�?�?   0  �   0 01090O0b0�0�0�0�0�0�0�0�0�0�0�0�0�033f4{4�4�4�4�4�4�485Q5i5�5�5�5�5�566*6<6E6^6s6{6�6�6�7�7�7�7	8"8;8S8l8�8�8�8�8�8�89K9]9o9x9�9�9�9�9:+:C:Y:o:�:�:�:�:;&;;;D;_;t;�;�;�;<)<D<n<�<�<�<�<�<�<�<==&=>=b>x>�>�>�>�>�>?%?>?Y?r?�?�?�?�?�?   @    0&0/0E0Q0_0x0�0�0�0�0�1�12-2E2^2w2�2�2�2�2�23#3I3Z3w3�3�3�3�3�3�3�34
4#424Z5p5�5�5�5�5�56666Q6j6�6�6�6�6�677&7<7N7V7o7�7�7�7�7�8�89$9<9U9n9�9�9�9�9�9::3:N:�:�:�:�:�:�:$;:;R;o;�;�;�;�;�;&<;<N<�<�<=#=A=W=i={=�=�=�=>>,>B>i>>�>�>�>�>??-???K?�?�?�?�?�?�?   P  $  0W0h0z0�0�0�0�011.1C1Y1o1�1�1�1�1�1�12]2u2�2�2�2�2�2�23C3Y3r3�3�3�3�3�34&4;4D4`4�4�4�4�4�4�405F5]5�5�5�5�5�5�5646K6�6�6�6�6�6�6�67K7]7o7x7�7�7�7�7818I8_8u8�8�8�8�8&9;9N9j99�9�9�9�9�9:#:+:D:Y:4;J;^;v;�;�;�;�;�;<<6<N<g<�<,=>=P=Y=n=�=�=�=�=�=
>>1>C>u>�>�>�>�>�>�>6?L?�?�?�? `  �   020v0�0�0�0�01�1�1�1�1�1�1�1=2S2l2�2�2�2�2�2�23343L3f3�3�3�3�344;4O4d4m4�4�4�4�4�4 5	5#5;5U5r5�5�5�5�5�5�56�6�6�6X7n7�7�7�78*8�8�8�8�8]9s9�9�9:=:a:�:�:H;�;�;<+<p<�<�<�<=<=^=m=�=�=�=>(>�>�>�>�>g?u?�?�?�?   p  t   0*0@0x0�0�0�01161L1�1�1�12#282C2w2�2�2�2�2�2$3=3f3�3&4r4�4&5Z5u5�5�5�5�5�5
6�6�6�6H7d7�7�7e<C=?d?�?�?�? �  �   0*0C0X0�0�01K1\1o1x1�1�1�1�1	2"272_2�2�2�2�2 3*3�3S4�4�4�4�5�5�517�78�8�8#9]9{9�9r:|:�:�;6<F<�<�<$=6=d=�=�=�=>%>>>U>g>y>�>? �  �   "0�01%1P1�1�1�12�2�2�2�263H3^3�4�4�4�4�465Z5�5 66}647v7�7�7�7�78&8P8�8�8?9�9&:8:N:`:r:�:�:;�;�;�;/<s< =F=X=n=�=�=�=�=)>�>�>?v? �  �   0F0X0�0�01'1?1�1�132�2�2�23/3E3Q6�6�6�6�6 777P7|7�7�78.8�8�8%9M9b9�9�9�9�9�9S::�:�:R;�;�<�<u=�=7>H>Z>s>�>�>a?�?�?�? �  �   �0�0h1}1�1�1�1�1�1�1F2_2w2�2�2�2�2
3373�3�3_4�5)8f8x8�8�8�8�8d9y9�9�9�9�9:4:M:e:~:�:�:�:�:;;0;E;�;�;�;�; <�<�<�<�<O=e=�=�=<>Z>�>�>�>-?�?�?   �  �   O00�0(1�1�1272�2383H3W3�3�3�3�34+4�4�4�4�4�4�4.5@5�5�5�5�5�506H6`6y6�6#787�7�78n8�8�8969b9�9�9":8:�:t;�;�;�;�;�;�;�;O<g<�<�<�<�<�<=�=�=�>�>z?�?�?�?�?�?�?�?   �  |   U0m0�0�0�0�01,1@1I1a1u1~1�1�12$2<2U2n2�2�2�2�2S3u344�5�5�5�5T67q7{7�7�7�7/8�8�8�8v9=;8<�<K=�=>�>?b?�?�?�?�?   �  �   M0f0�0�0&1>1\1�1�1<2W2k2t2�2�2�23)3A3Z3�3�3�3�3�3�3N4f44�4�4O5d5x5�5�5�5�5�516M6a6z6�697s7�7�8�8�8�89949f9t9�9�9�9�9�9:�;�;�;�;k<�<�<�<�<�<�<=I>T>�>�>	??1?D?�?�?�?�? �  @   �0�2�234(4e5�536p67C7J7|7�7�7~9�9F:X:r:�>?"?4?B?l?     4   �3�4�4e577�78�8�8�8�9�9h:�:;%;�;�;�?�?    ,   v3�3w7�78%8q8�8�8�8�8v9�9U:V;e;�?     x   b0�1�1�12V2e2x2�2�2�2�2�23373?3E3J3[3�3�3�3F4Z4�466�6�6717<7K7k7v7�7�7�7�7�78Q8�89F9U9l9�9�9:;;�=�=   0 p   f1x1�1�1�1�1�1�1�1-2:2N2�23�3�34414P4�4�5�5�6�6]7&8589�9&:8:x;==�=�=�= >>u>�>�>�>�>�> ??�?�?�?   @ `   *1V1h1�2�45v8�8v:�:V;f;$<A<M<W<�<�<�<�<�<7=M=\=�=�=�=>$>�>�>�>�>�>�>�>?4?J?q?�?�?�?   P �   090d0�0�0�0�01$1D1d1�1�1�1�1242d2�2�2�2D3�3�3�3�3�3D4Y4y4�4�4545T5�5�5�56$6D6d6�6�6�6�67D7t7�7�7�7848d8�8�8�89$9T9�92:f:L;x;�;==%=H=R=q=�=�=�=>D>�>�>$?K?�?�?�?   ` \   0+0T0|0�01T1�1�12�23�34�5�5*6�6�657�7�7;8{8�8�89[9�9�9I:�:�:;h;�=>>>?a?   p p   �01A1z1�1�2�203s3�34c4�4#5�5�5#6�6�6C7�78c8�8#9�9�93:�:�:Y;�;�;i<�<=@=z=�=�= >0>d>�>�>?A?{?�?�?�?   � �   .0j0�0�0;1�1�12^2�2�2343q3�3�34T4�4�4&5T5�5%6*656K6h6r6�6 8�8�8�8�8�8�8�8�8�8�8&9�98:<:@:D:H:L:P:T:X:�:;";D;o;�;�;�;�;<!<A<d<�<�<�<=4=d=�=�=>4>a>�>�>�>t?�?�?�?   � �   040d0�0�0�011*1H1a1s1�1�1�1�1�122=2V2h2|2�2�2�23T3�3�3�3�344�4�45D5\5�5�56D6q6�6�6t7�78�8�9X:�:�:�:�:�:�:9;�;�;�;�;
<<D<d<�<(=�=	>4>d>�>�>�>:?T?   � �   �01D1�1�1�1�1�1\2a3�3�3�3�3�34#434�4�4�4�455'595P5�5�5�5�5 66_6x6�6.7B7T7e7�7�7�78/8?8f8�8�8�8f9�9�<�<�<=C=m=�=�=�?�?�?�? � p   0080W0�0�0�0�0�0�011/1A1S1b1u154:M:v:�:�:�:�:�::;o;�;�;�;<<_<q<�<�<�<�<(=;=|>�>�>�>+?G?�?�?�?�?   � �   040E0d0u0�0�0�0�0�01D1q1�1�1�1�1�12!242T2t2�2�2�2�2	343d3�3�3�34!444T4�4�4�4�4545d5�5�5�5�5646T6t6�6�6�6�6747T7w7�7�7�7�78888�8�8�89%9d9�9�9�9�9$:A:[:T;t;�;�;�;�;<4<T<�<�<�<=$=D=t=�=�=�=>!>D>d>�>�>�>�>?$?D?d?�?�?�?�?   � �   00+0H0�0�0�0151t1�1�1�1�142Q2k2d3�3�3�3�34$4D4d4�4�4�4�455/5=5L5t5�5�5�5�5�56A6a6�6�6�6�6�6�6747T7i7�7�7�7�7�7848T8t8�8�8�8�8949T9g9}9�9�9�9�9�9:4:R:f:v:�:�:;1;Q;t;�;�;�;�;<4<T<t<�<�<�<�<=4=T=t=�=�=�=><>d>�>�>�>�>?4?T?t?�?�?�?   � �   040T0t0�0�0�0�0$1D1d1�1�1�1�1212T2�2�2�2�23$3F3Z3j3�3�3�3�3�34)4@4O4�4�4�45D5o5�5�5�567.7<7T7q7�7�7�7$8T88�8�89D9h9�9�:�:�:�:�:�:;o;�;�;�;<<1<M<x<�<�<�<�<=/=\=�=�=�=3>E>�>�>)?E?�?�?   � �   )0L0h0�0�0�0�01m1�12\2�2�23$3D3d3�3�3�3�34$4D4a4t4�4�4�4545O5o5�5�5�5�56B6d6�6�6�6�67$7D7t7�7�7�7848t8�8�8�8949T9t9�9�9�9�9:1:D:d:�:�:�:.;N;c;�;<a<�<�<X=z=�=>:>]>�>�>?~?�?�?     �   30\0y0�0�01�1�1�1S2|2�23<3Y3�3�34{4�45q5�5�56q6�6�6\7�7�78�8�8�8>9^9s9�9!:�:�:$;D;a;q;�;�;�;�;<4<d<�<�<�<=$=D=a=�=�=�=C>`>�>�>�>�>	?F?U?�?�?�?�?  �   040T0�0�0�0�01A1d1�1�1�1�12$2T2t2�2�23$3D3a3q3�3�3�3(4g4�4�45D5a5t5�5�5�5616T6t6�6�6�6$7T7�7�7�7�7848T8t8�8�8�8�89919A9T9t9�9�9�9:!:4:t:�:�:�:�:;;$;D;d;�;�;�;�;<4<T<t<�<�<�<�<=/=Q=d=�=�=�=>4>T>t>�>�>�>�>?4?T?t?�?�?�?   �   0T0�0�01T1�1�1�12A2a2t2�2�2�2�23$3D3d3�3�3�3�3B4h4�4�4�4�45T5t5�5�5�5�566&6T6t6�6�6�67/7G7[7k7�7�7�78*8H8]8�8�8�8�8�8�89"9D9�9�9�9+:=:Q:a:�:�:�:;!;1;d;�;�;�;C<U<�<�<�<�<=4=T=t=�=�=�=�=>!>4>t>�>�>�>�>?Y?�?�?�?�? 0 �   0!010D0a0t0�0�0�0�011(1A12B2r2�2�2"3U3�3�3%454u4�45M5�5�56R6�6�67E7�7�78R8�8�8�829e9�9�95:u:�:�:8;S;�;�;�;�;<U<�<�<=e=�=�=A>i>�>�>�>�>�>?<?d?�?�?�?   @ �   	0H0o0�0�01U1}1�1�12B2v2�2�2u3�3�3�3�34$4D4d4�4�4�4�4�4�45545X5q5�5�5�5�56D6d6�6�6�6�67$7d7�7�7�7�7�788A8_8�8�8�8�8949T9�9�9�9�9�9:%:L:\::�:�:�:�:;&;T;j;�;�;�;< <q<�<�<�<�<==C=c=w=�=�=�=�=>4>T>�>�>�>?4?T?�?�?�?�?   P �   0$0d0�0�0$1d1�1�1�1�12$2D2d2�2�2�2343T3�3�3�3�3!4D44�4�4�45W5�5�5�56T6�6�6�6717T7q7�7�7�7�7848d8�8�8�8B9a9�9�9�9�9:A:a:�:�:�:�:;D;t;�;�;�;<&<a<�<�<$=Q=t=�=�=�=!>A>q>�>�>�>?!?D?�?�?�?�? ` �   $0T0t0�0�01A1a1�1�1�12$22272T2}2�2�2$3T3t3�3�34W4�4W5�5�5�5�5646]6�6�6�6$7A7d7�8�89$9T9�9�9�9�9:4:T:u:�:�:�:;4;Q;t;�;�;<1<T<�<�<�<�<!=4=T=�=�=D>�>�>�>�>?4?{?�? p �   0.0X0s0�0�0�011<1V1�1�1�1�1
22O2c2x2�2�233;3U3r3�3�3[4l4�4�4�4�45m5l7�9�9�9�91:A:x:�:�:,<0<4<8<k<p<�<�<�<=4=T=t=�=�=�=�=>:>�>�>Z?�? � �   0T0�0�0�01!1D1d1�1�1�1�1242T2t2�2�2�2313�3�314X4�4(5�5�5,6G6�67d7�7�7-8A8Q8m8�8�8;�;�;�;<K<�<�<�<�<�<�<=!=.=F=Y=k=}=�=�=�=�=�= >>2>D>V>t>�>�>�>�>�>�>�>�>?1?C?`?x?�?�?�?�?�?�? �   0%0<0V0h0{0�0�0�0�0�0�011(1E1a1s1�1�1�1�1�1�1
2'282U2l2�2�2�2�2�2�2�2323]3�3�3�3�3�3�3�3�34%4A4S4p4�4�4�4�4�4�45555L5f5x5�5�5�5�5�5�5606=6Y6z6�6�6�67!7�7�7�7�7�7�7�78!8*8=8�8�8�8�89�9�9 :Q:�:�:�:�:�:!;4;T;q;�;�;�;�;T<B=I=P=W=^=e=l=s=�=�=�=�>)?�?�?   � x   0!0O0q0�0191�12�2�2�2�2�2�2�23<3l3�3�3�3�324N4X4f4k4�4�4�4595a5�5�5�5�52686d6q6w6�6�6�6�67%7?7X7\7`7d7h7l7 � ,   �1�13]4d4�4�4g5q5�5�5�5�5?1?]?�?�? � d   0e0�0�0"1R1�1�1252u2�2�223b3�3�3�354u4�45U5�5�56U6�67�;<< <$<(<�=�=�=�=!?4?a?�?�?�?�? � �   030F0q0�0�0�01$1T1�1�1�1�1$2T2�2�2�2�2$3d3�3�3�3�34$4D4t4�4�4�4a5t5�5�566�7�7808�9�:;b;�;�<�<�<S=k=�=�=!>+>�>�>�>d?�?�?�? � �   �3]4m4�5�556d6k6�6�6�6�6-7}7B9J9T9c9p9v9�9�9�9�9Y:d:u:�:�:�:�:�:;';@;H;`;q;�;�;�;�;�;<I<S<g<�<�<�<�<=+=�=�=Q?^?q?�?�?�?�?�?�? � �   0U0e0}0�0�0:1J1Z1j1v1�1�1�1�1�1�1�2O3g3l3�5�5.6@6�6�6�6�6<79�9L:Q:W:[:a:e:k:o:u:y:~:�:�:�:�:�:�:�:�:�:�:/;H;O;W;\;`;d;�;�;�;�;�;�;�;�;�;�;�;><D<H<L<P<�<�<�<�<�<�<�<=;=m=t=x=|=�=�=�=�=�=�=�=�=�=�=A>U>�>�>?,?I?V?�?   `   C1U1'212>2Y2`2x2�2�2�23W3]3n3�3�3�34!4�4�4�45%5�5�5�5�6�7�7�7�7G8�8�8�9=;�<�=;?E?�?    �   ;0@0J0~0�0�0�0�0�01;1W1o1�1�1b2�2�2G3a3j3r3�3�3>4P4�4�4�4�45J66�6�6�6�6�6�6�67!7(7,7074787<7@7D7�7�7�7�7�788,83888<8@8a8�8�8�8�8�8�8�8�8�8�8*9094989<9�9�9�9?:X:�:�:�:�:�:;p;�;�;�;�;�;<<<(<0<;<k<�<2=�=>�>T?�?�?   �   U0a0�0�0S1_1�1�1X2d2�2j35�5�5�56-656S6[6�6�6�6�6�6�6!7*767s7|7�778B8e8)969K9]9{9�9�9�:�:2;~;�;<�<�<�<=,=5=>=J=V=b=n=y=&>�>?A?�?�?�?�?   0 L   0-0>0�0�0_1`23�4$5k5�5�56�6�6�6�6%8�8�899#9,9�9:;';�;>>1>�> @ �   01a1�2|4�7�7�7�9�:�:�:�:�:�:;;:;@;K;W;l;s;�;�;�;�;�;�;�;�;�;�;�;<<<!<+<2<J<Y<`<m<�<�<�<==;=A=]=u=�=>8>B>z>�>�>�>�>�>�>??!?/?:?A?\?a?i?o?v?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   P �   	000$0)04090F0T0Z0g0�0�0�0�011G1R1�1�1�1�1�1�1�1�1�1�1�1 22222+24292?2I2R2]2i2n2~2�2�2�2�2�2�2�2�24W4n4�5�5,696C6Q6Z6d6�6�6�6�6�6�67>7s7�7�78[8�8�8[9g9z9�9�9�9�9�9�9:::: :/:V::�:�:�:;;e<=�? ` �   0K0�5`68R8[8�8�8�8�8:8:=:K:S:_:f:o:�:�:�:�:�:�:�:�:�:�:�:;;;>;E;^;r;x;�;�;�;M<m<{<�<�>�>�>�>�>???&?8?K?V?\?b?g?p?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   p �   00030D0J0[0�0\4h4�4�4�4@577&797V7�7�8�8�8�89-939M9\9i9u9�9�9�9�9�9�9�9�9::=:p::�:�:�:�;�;<#<D<J<|<�<�<=%=M=f=�=�=�=;>A>e>�>�>�?�? � P   K0�01�1�1�2�2H3�4�56�6�67&7�7�7&8�8�8�8*949�9:�:�;�<u=�=�=�=�=>?�? � $   �041q1{1�1�1�12\3�3�3!4;   � �   O5V5u5~5�5�5�5�5�5�5]6e6x6�6�6�6�6�6�6�6�6�6�677717q7~7�7�7�7�7�7g8t8|8�8�8�89(929C9N9;;; ;%;+;�;�;�;�;�;�;�;�;,<{<�<�<�<�<�<==K=�=�=�=�=�>�>�>�>�>??5?=?v?~?�?�? � �   (0X0a0|0�0�0�0�0�0�0�0
1%1,151>1G1P1Y1e1q1z1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�122}2�2-3E3P3t3}3�3�3�3�3�34D4W4o4�4�4�4�4�5N6l6�6�67 7k:[;�<=9=? � T   11 1$1(1,10141D1�1u2�2�2�23D3J3�3�3<4�4�4�4�4556�6(7�7�7.868E8M8�8�8�? � �   )1D1�162@2b2�2�3�3M4�4�45�5�6�677%767E7b7�7�7�7�8�8�9::":,:4:A:H:x:;�;�;L<a<�<�<�<=A=y=�=�=;>A>e>�>�>�>�>?�?�?�?�?�?�?   � \   0M0R0�0�0�0�0�0�0#1,121s7�7�7�78J8^9i9r9�9�9:!:3:E:W:i:�:�<�< =&?<?M?j?�?�?�?�?   � 4   =0|0�0�0I1n13Z344^4g4�4�4;5D5]5�5�5�5�51;   X   g<k<o<s<w<{<<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<9=�>0?O?n?�?�?    d   	00J0Z0�0�0�0�0�0�011=1I2�2=3I3�3�3�3�5�5_6�8�:�:�:�:�;�;�;�;�;�;P<q<}<�<�<�<�<,=b=�>�?�?     �   a0p0�0�0�1�1t2�2�23�3�3434q4�4n5�5�5�5�5�5�56
66*61676M6h67{7�7�7�7�778G8b8�8�8�8$9@9�9�9�9�9�9+:=:�:�:�:;;L;n<? 0 �   k0�0�0�0�0%1.2�2�243�3�5�5�5�5�5�5(6b6p6v6�6�6�6�6�6�6�6�6�6�6�6�677V7s7�7�7�7�78879U9�9�9�9�9:::#:�:�:m;a<�=�>   @ L   �1V2�2�2�233'3g3�3j6�6�6�6
77,7Q7h78F9B:;<<�<�=J>P>�>�>?�?�? P P   b0X1`12�2�3�364<4L4�4535�5�8�8�;�;�;�;<<
<<<<<<+<==-=Y=�=�=   ` 0   �7�9�9�9�9�9�9�:�:;&;�;�;�;�<�=�=�?�?   p L   %0S0�0�0�0�1�1�1222�2�2�2!3]3�3�3�34�4+5�5�6Q9�:�;r<�>3?k?�?�?   � l   (0�0�0Y1�12d2�293�4&5l6�78[8�8�8�89:9s9�9:D:t:�:�:$;J;z;�;<@<j<�<�<�<;=s=�=�=�=*>u>�>�>?i?�?�? � H   0=0r0�0�0�0�0#1F1i1�1�1�1222'232?2I2U2b2j2t2�2�2�2�2�2�2�2   � �  `1d1h1l1p1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 286<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888�8�8�:�:�:�:�:�:�:�:�:@;D;H;L;P;T;X;\;`;d;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<< <$<(<,<0<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<h=l=p=t=x=�=�=�=�=�=�=�=�=�=�=�=�=X>\>x>|>�>�>�>�?�?�?�?�?�?�?�?�?�? � T    000�0�0�0�0�0�0�0�0�0�0 1�9�9�9�9�9�9�9�9�9�9�9 ::::::�:�:�:�:4;8;   � �   �9�9�9�9�9�9�9 :::: :(:0:8:@:H:P:X:`:h:p:x:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;; ;(;0;8;@;H;P;X;`;h;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�< � �  �2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�5�5�6�6�6�6�6�6�6�6�6�6�67777 7(7@7D7\7l7p7�7�7�7�7�7�7�7�7�7�7�78888,8<8@8P8T8X8`8x8|8�8�8�8�8�8�8�8�8�8�8�8�899 989H9L9P9T9\9t9x9�9�9�9�9�9�9�9�9�9�9�9�9: :$:4:8:@:X:h:l:|:�:�:�:�:�:�:�:�:�:�:�:�:;;;; ;$;(;,;4;L;\;`;p;t;x;�;�;�;�;�;�;�;�;�;�;�;<<<<0<@<D<T<X<\<`<h<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ====(=8=<=@=H=`=d=|=�=�=�=�=�=�=�=�=�=�=�=�=>>> >$>,>D>T>X>h>l>t>�>�>�>�>�>�>�>�>�>�>�> ????(?8?<?D?\?l?p?�?�?�?�?�?�?�?�?�?�?�? � �   00000$0<0L0P0`0d0t0x0�0�0�0�0�0�0�0�0�0�0111(181<1L1P1T1\1t1�1�1�1�1�1�1�1�1�1�1�1�1222,2024282@2X2h2l2|2�2�2�2�2�2�2�2�2�2�2�2 333$3(3,343L3�4�4�455$5H5h5p5x5�5�5�5�5�5�5�5�5�5�5�5�5�56666$6,646<6D6L6T6\6d6l6t6|6�6�6�6�6�6�6�6�6�6�6�677$7,747<7D7L7T7\7d7p7�7�7�7�7�7�7�7 88848<8H8h8p8x8�8�8�8�8�8 9 9(90989@9H9P9X9`9h9p9x9�9�9�9�9�9�9�9�9�9�9�9:: :(:0:8:@:H:T:t:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;$;,;4;<;D;P;p;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<8<@<H<P<X<`<h<p<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ==== =(=0=8=@=H=P=X=`=h=p=x=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>$>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�> ???? ?(?0?8?@?H?P?X?`?h?p?x?�?�?�?�?�?�?�?�?�?�?�?�?�?   � �  0000$0,040<0D0L0T0\0h0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�233(3L3l3t3|3�3�3�3�3�3�3�3�3�3�3�3�3 44444<4D4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4�4�4�45$5,545<5D5L5T5\5d5l5x5�5�5�5�5�5�5�5666 6(606<6\6d6l6t6|6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�780888@8H8P8X8`8h8p8x8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99949<9D9L9T9\9d9l9t9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9::::$:0:P:X:`:h:t:�:�:�:�:�:�:�:�:�:�:; ;H;X;�;�;�;�;�;�;�;<<,<8<`<t<�<�<�<�<�<�<�<�<�<=(=0=8=@=H=P=\=|=�=�=�=�=�=�=�=>><>D>L>P>T>\>p>x>�>�>�>�>�>�>�>�> ???$?,?4?@?h?|?�?�?�?�?�?�?�?�?�?   �  00000080L0T0`0�0�0�0�0�0�01$1H1\1l1|1�1�1�1�1�1�122,2@2H2`2l2�2�2�2�2�2�23,343D3X3`3�3�3�3�3�3�3�34,484X4h4t4�4�4�4�4�45(545<5T5\5�5�5�5�5�5�56 6(646T6\6h6�6�6�6�6�6�6�6�67$707P7\7|7�7�7�7�7�7�7�788 8$8(808D8`8�8�8�8�8�89(9H9h9�9�9�9�9�9:(:4:@:`:�:�:�:�:�:�:�:�:�: ;(;,;D;H;d;h;p;x;�;�;�;�;�;�;�;�;<<,<0<P<p<�<�<�<�<�<�<=0=P=p=�=�=�=�=>0>P>p>�>�>�>�>�>�>?0?P?\?t?x?�?   (   00 080<0@0\0x0�0�0�0�01L1�1�1�102P2�2�2 3 3@3d3�3�3�3�3�3�34 4$4(4D4`4x4�4�4�4�4�4�4�4�4�4�4�4�4�45585<5@5D5H5L5P5T5X5p5t5x5|5�5�5�5�5�5�5�566686@6D6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�677P7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88<�=�=�=�=�=�=>>>>> >$>�?�?�?�?�?�?�?�?�?�? 0 l  �0�0�3�3�3�3�3�3�3�34444$4,444<4D4L4T4\4d4l4t4|4�4�45"5&5*5.52565:5>5B5F5J5N5R5V5Z5^5b5f5j5n5r5v5z5~5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�566
66666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 777L8T8\8d8l8t8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�89999$9,9::                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    